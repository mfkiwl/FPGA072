
module gbuf (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
