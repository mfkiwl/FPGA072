// Copyright (C) 2018  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details.

// VENDOR "Altera"
// PROGRAM "Quartus Prime"
// VERSION "Version 18.1.0 Build 625 09/12/2018 SJ Standard Edition"

// DATE "05/22/2020 12:53:10"

// 
// Device: Altera 5AGXMA7G4F31C4 Package FBGA896
// 

// 
// This greybox netlist file is for third party Synthesis Tools
// for timing and resource estimation only.
// 


module nco_test (
	clk,
	clken,
	phi_inc_i,
	fsin_o,
	fcos_o,
	out_valid,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	clk;
input 	clken;
input 	[31:0] phi_inc_i;
output 	[17:0] fsin_o;
output 	[17:0] fcos_o;
output 	out_valid;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \nco_ii_0|dop|sin_o[0]~q ;
wire \nco_ii_0|dop|sin_o[1]~q ;
wire \nco_ii_0|dop|sin_o[2]~q ;
wire \nco_ii_0|dop|sin_o[3]~q ;
wire \nco_ii_0|dop|sin_o[4]~q ;
wire \nco_ii_0|dop|sin_o[5]~q ;
wire \nco_ii_0|dop|sin_o[6]~q ;
wire \nco_ii_0|dop|sin_o[7]~q ;
wire \nco_ii_0|dop|sin_o[8]~q ;
wire \nco_ii_0|dop|sin_o[9]~q ;
wire \nco_ii_0|dop|sin_o[10]~q ;
wire \nco_ii_0|dop|sin_o[11]~q ;
wire \nco_ii_0|dop|sin_o[12]~q ;
wire \nco_ii_0|dop|sin_o[13]~q ;
wire \nco_ii_0|dop|sin_o[14]~q ;
wire \nco_ii_0|dop|sin_o[15]~q ;
wire \nco_ii_0|dop|sin_o[16]~q ;
wire \nco_ii_0|dop|sin_o[17]~q ;
wire \nco_ii_0|dop|cos_o[0]~q ;
wire \nco_ii_0|dop|cos_o[1]~q ;
wire \nco_ii_0|dop|cos_o[2]~q ;
wire \nco_ii_0|dop|cos_o[3]~q ;
wire \nco_ii_0|dop|cos_o[4]~q ;
wire \nco_ii_0|dop|cos_o[5]~q ;
wire \nco_ii_0|dop|cos_o[6]~q ;
wire \nco_ii_0|dop|cos_o[7]~q ;
wire \nco_ii_0|dop|cos_o[8]~q ;
wire \nco_ii_0|dop|cos_o[9]~q ;
wire \nco_ii_0|dop|cos_o[10]~q ;
wire \nco_ii_0|dop|cos_o[11]~q ;
wire \nco_ii_0|dop|cos_o[12]~q ;
wire \nco_ii_0|dop|cos_o[13]~q ;
wire \nco_ii_0|dop|cos_o[14]~q ;
wire \nco_ii_0|dop|cos_o[15]~q ;
wire \nco_ii_0|dop|cos_o[16]~q ;
wire \nco_ii_0|dop|cos_o[17]~q ;
wire \nco_ii_0|ux710isdr|data_ready~q ;
wire \clk~input_o ;
wire \reset_n~input_o ;
wire \clken~input_o ;
wire \phi_inc_i[31]~input_o ;
wire \phi_inc_i[30]~input_o ;
wire \phi_inc_i[29]~input_o ;
wire \phi_inc_i[28]~input_o ;
wire \phi_inc_i[27]~input_o ;
wire \phi_inc_i[26]~input_o ;
wire \phi_inc_i[25]~input_o ;
wire \phi_inc_i[24]~input_o ;
wire \phi_inc_i[23]~input_o ;
wire \phi_inc_i[22]~input_o ;
wire \phi_inc_i[21]~input_o ;
wire \phi_inc_i[20]~input_o ;
wire \phi_inc_i[19]~input_o ;
wire \phi_inc_i[18]~input_o ;
wire \phi_inc_i[17]~input_o ;
wire \phi_inc_i[16]~input_o ;
wire \phi_inc_i[15]~input_o ;
wire \phi_inc_i[14]~input_o ;
wire \phi_inc_i[13]~input_o ;
wire \phi_inc_i[12]~input_o ;
wire \phi_inc_i[11]~input_o ;
wire \phi_inc_i[10]~input_o ;
wire \phi_inc_i[9]~input_o ;
wire \phi_inc_i[8]~input_o ;
wire \phi_inc_i[7]~input_o ;
wire \phi_inc_i[6]~input_o ;
wire \phi_inc_i[5]~input_o ;
wire \phi_inc_i[4]~input_o ;
wire \phi_inc_i[3]~input_o ;
wire \phi_inc_i[2]~input_o ;
wire \phi_inc_i[1]~input_o ;
wire \phi_inc_i[0]~input_o ;


nco_test_nco_test_nco_ii_0 nco_ii_0(
	.sin_o_0(\nco_ii_0|dop|sin_o[0]~q ),
	.sin_o_1(\nco_ii_0|dop|sin_o[1]~q ),
	.sin_o_2(\nco_ii_0|dop|sin_o[2]~q ),
	.sin_o_3(\nco_ii_0|dop|sin_o[3]~q ),
	.sin_o_4(\nco_ii_0|dop|sin_o[4]~q ),
	.sin_o_5(\nco_ii_0|dop|sin_o[5]~q ),
	.sin_o_6(\nco_ii_0|dop|sin_o[6]~q ),
	.sin_o_7(\nco_ii_0|dop|sin_o[7]~q ),
	.sin_o_8(\nco_ii_0|dop|sin_o[8]~q ),
	.sin_o_9(\nco_ii_0|dop|sin_o[9]~q ),
	.sin_o_10(\nco_ii_0|dop|sin_o[10]~q ),
	.sin_o_11(\nco_ii_0|dop|sin_o[11]~q ),
	.sin_o_12(\nco_ii_0|dop|sin_o[12]~q ),
	.sin_o_13(\nco_ii_0|dop|sin_o[13]~q ),
	.sin_o_14(\nco_ii_0|dop|sin_o[14]~q ),
	.sin_o_15(\nco_ii_0|dop|sin_o[15]~q ),
	.sin_o_16(\nco_ii_0|dop|sin_o[16]~q ),
	.sin_o_17(\nco_ii_0|dop|sin_o[17]~q ),
	.cos_o_0(\nco_ii_0|dop|cos_o[0]~q ),
	.cos_o_1(\nco_ii_0|dop|cos_o[1]~q ),
	.cos_o_2(\nco_ii_0|dop|cos_o[2]~q ),
	.cos_o_3(\nco_ii_0|dop|cos_o[3]~q ),
	.cos_o_4(\nco_ii_0|dop|cos_o[4]~q ),
	.cos_o_5(\nco_ii_0|dop|cos_o[5]~q ),
	.cos_o_6(\nco_ii_0|dop|cos_o[6]~q ),
	.cos_o_7(\nco_ii_0|dop|cos_o[7]~q ),
	.cos_o_8(\nco_ii_0|dop|cos_o[8]~q ),
	.cos_o_9(\nco_ii_0|dop|cos_o[9]~q ),
	.cos_o_10(\nco_ii_0|dop|cos_o[10]~q ),
	.cos_o_11(\nco_ii_0|dop|cos_o[11]~q ),
	.cos_o_12(\nco_ii_0|dop|cos_o[12]~q ),
	.cos_o_13(\nco_ii_0|dop|cos_o[13]~q ),
	.cos_o_14(\nco_ii_0|dop|cos_o[14]~q ),
	.cos_o_15(\nco_ii_0|dop|cos_o[15]~q ),
	.cos_o_16(\nco_ii_0|dop|cos_o[16]~q ),
	.cos_o_17(\nco_ii_0|dop|cos_o[17]~q ),
	.data_ready(\nco_ii_0|ux710isdr|data_ready~q ),
	.clk(\clk~input_o ),
	.reset_n(\reset_n~input_o ),
	.clken(\clken~input_o ),
	.phi_inc_i_31(\phi_inc_i[31]~input_o ),
	.phi_inc_i_30(\phi_inc_i[30]~input_o ),
	.phi_inc_i_29(\phi_inc_i[29]~input_o ),
	.phi_inc_i_28(\phi_inc_i[28]~input_o ),
	.phi_inc_i_27(\phi_inc_i[27]~input_o ),
	.phi_inc_i_26(\phi_inc_i[26]~input_o ),
	.phi_inc_i_25(\phi_inc_i[25]~input_o ),
	.phi_inc_i_24(\phi_inc_i[24]~input_o ),
	.phi_inc_i_23(\phi_inc_i[23]~input_o ),
	.phi_inc_i_22(\phi_inc_i[22]~input_o ),
	.phi_inc_i_21(\phi_inc_i[21]~input_o ),
	.phi_inc_i_20(\phi_inc_i[20]~input_o ),
	.phi_inc_i_19(\phi_inc_i[19]~input_o ),
	.phi_inc_i_18(\phi_inc_i[18]~input_o ),
	.phi_inc_i_17(\phi_inc_i[17]~input_o ),
	.phi_inc_i_16(\phi_inc_i[16]~input_o ),
	.phi_inc_i_15(\phi_inc_i[15]~input_o ),
	.phi_inc_i_14(\phi_inc_i[14]~input_o ),
	.phi_inc_i_13(\phi_inc_i[13]~input_o ),
	.phi_inc_i_12(\phi_inc_i[12]~input_o ),
	.phi_inc_i_11(\phi_inc_i[11]~input_o ),
	.phi_inc_i_10(\phi_inc_i[10]~input_o ),
	.phi_inc_i_9(\phi_inc_i[9]~input_o ),
	.phi_inc_i_8(\phi_inc_i[8]~input_o ),
	.phi_inc_i_7(\phi_inc_i[7]~input_o ),
	.phi_inc_i_6(\phi_inc_i[6]~input_o ),
	.phi_inc_i_5(\phi_inc_i[5]~input_o ),
	.phi_inc_i_4(\phi_inc_i[4]~input_o ),
	.phi_inc_i_3(\phi_inc_i[3]~input_o ),
	.phi_inc_i_2(\phi_inc_i[2]~input_o ),
	.phi_inc_i_1(\phi_inc_i[1]~input_o ),
	.phi_inc_i_0(\phi_inc_i[0]~input_o ));

assign \clk~input_o  = clk;

assign \reset_n~input_o  = reset_n;

assign \clken~input_o  = clken;

assign \phi_inc_i[31]~input_o  = phi_inc_i[31];

assign \phi_inc_i[30]~input_o  = phi_inc_i[30];

assign \phi_inc_i[29]~input_o  = phi_inc_i[29];

assign \phi_inc_i[28]~input_o  = phi_inc_i[28];

assign \phi_inc_i[27]~input_o  = phi_inc_i[27];

assign \phi_inc_i[26]~input_o  = phi_inc_i[26];

assign \phi_inc_i[25]~input_o  = phi_inc_i[25];

assign \phi_inc_i[24]~input_o  = phi_inc_i[24];

assign \phi_inc_i[23]~input_o  = phi_inc_i[23];

assign \phi_inc_i[22]~input_o  = phi_inc_i[22];

assign \phi_inc_i[21]~input_o  = phi_inc_i[21];

assign \phi_inc_i[20]~input_o  = phi_inc_i[20];

assign \phi_inc_i[19]~input_o  = phi_inc_i[19];

assign \phi_inc_i[18]~input_o  = phi_inc_i[18];

assign \phi_inc_i[17]~input_o  = phi_inc_i[17];

assign \phi_inc_i[16]~input_o  = phi_inc_i[16];

assign \phi_inc_i[15]~input_o  = phi_inc_i[15];

assign \phi_inc_i[14]~input_o  = phi_inc_i[14];

assign \phi_inc_i[13]~input_o  = phi_inc_i[13];

assign \phi_inc_i[12]~input_o  = phi_inc_i[12];

assign \phi_inc_i[11]~input_o  = phi_inc_i[11];

assign \phi_inc_i[10]~input_o  = phi_inc_i[10];

assign \phi_inc_i[9]~input_o  = phi_inc_i[9];

assign \phi_inc_i[8]~input_o  = phi_inc_i[8];

assign \phi_inc_i[7]~input_o  = phi_inc_i[7];

assign \phi_inc_i[6]~input_o  = phi_inc_i[6];

assign \phi_inc_i[5]~input_o  = phi_inc_i[5];

assign \phi_inc_i[4]~input_o  = phi_inc_i[4];

assign \phi_inc_i[3]~input_o  = phi_inc_i[3];

assign \phi_inc_i[2]~input_o  = phi_inc_i[2];

assign \phi_inc_i[1]~input_o  = phi_inc_i[1];

assign \phi_inc_i[0]~input_o  = phi_inc_i[0];

assign fsin_o[0] = \nco_ii_0|dop|sin_o[0]~q ;

assign fsin_o[1] = \nco_ii_0|dop|sin_o[1]~q ;

assign fsin_o[2] = \nco_ii_0|dop|sin_o[2]~q ;

assign fsin_o[3] = \nco_ii_0|dop|sin_o[3]~q ;

assign fsin_o[4] = \nco_ii_0|dop|sin_o[4]~q ;

assign fsin_o[5] = \nco_ii_0|dop|sin_o[5]~q ;

assign fsin_o[6] = \nco_ii_0|dop|sin_o[6]~q ;

assign fsin_o[7] = \nco_ii_0|dop|sin_o[7]~q ;

assign fsin_o[8] = \nco_ii_0|dop|sin_o[8]~q ;

assign fsin_o[9] = \nco_ii_0|dop|sin_o[9]~q ;

assign fsin_o[10] = \nco_ii_0|dop|sin_o[10]~q ;

assign fsin_o[11] = \nco_ii_0|dop|sin_o[11]~q ;

assign fsin_o[12] = \nco_ii_0|dop|sin_o[12]~q ;

assign fsin_o[13] = \nco_ii_0|dop|sin_o[13]~q ;

assign fsin_o[14] = \nco_ii_0|dop|sin_o[14]~q ;

assign fsin_o[15] = \nco_ii_0|dop|sin_o[15]~q ;

assign fsin_o[16] = \nco_ii_0|dop|sin_o[16]~q ;

assign fsin_o[17] = \nco_ii_0|dop|sin_o[17]~q ;

assign fcos_o[0] = \nco_ii_0|dop|cos_o[0]~q ;

assign fcos_o[1] = \nco_ii_0|dop|cos_o[1]~q ;

assign fcos_o[2] = \nco_ii_0|dop|cos_o[2]~q ;

assign fcos_o[3] = \nco_ii_0|dop|cos_o[3]~q ;

assign fcos_o[4] = \nco_ii_0|dop|cos_o[4]~q ;

assign fcos_o[5] = \nco_ii_0|dop|cos_o[5]~q ;

assign fcos_o[6] = \nco_ii_0|dop|cos_o[6]~q ;

assign fcos_o[7] = \nco_ii_0|dop|cos_o[7]~q ;

assign fcos_o[8] = \nco_ii_0|dop|cos_o[8]~q ;

assign fcos_o[9] = \nco_ii_0|dop|cos_o[9]~q ;

assign fcos_o[10] = \nco_ii_0|dop|cos_o[10]~q ;

assign fcos_o[11] = \nco_ii_0|dop|cos_o[11]~q ;

assign fcos_o[12] = \nco_ii_0|dop|cos_o[12]~q ;

assign fcos_o[13] = \nco_ii_0|dop|cos_o[13]~q ;

assign fcos_o[14] = \nco_ii_0|dop|cos_o[14]~q ;

assign fcos_o[15] = \nco_ii_0|dop|cos_o[15]~q ;

assign fcos_o[16] = \nco_ii_0|dop|cos_o[16]~q ;

assign fcos_o[17] = \nco_ii_0|dop|cos_o[17]~q ;

assign out_valid = \nco_ii_0|ux710isdr|data_ready~q ;

endmodule

module nco_test_nco_test_nco_ii_0 (
	sin_o_0,
	sin_o_1,
	sin_o_2,
	sin_o_3,
	sin_o_4,
	sin_o_5,
	sin_o_6,
	sin_o_7,
	sin_o_8,
	sin_o_9,
	sin_o_10,
	sin_o_11,
	sin_o_12,
	sin_o_13,
	sin_o_14,
	sin_o_15,
	sin_o_16,
	sin_o_17,
	cos_o_0,
	cos_o_1,
	cos_o_2,
	cos_o_3,
	cos_o_4,
	cos_o_5,
	cos_o_6,
	cos_o_7,
	cos_o_8,
	cos_o_9,
	cos_o_10,
	cos_o_11,
	cos_o_12,
	cos_o_13,
	cos_o_14,
	cos_o_15,
	cos_o_16,
	cos_o_17,
	data_ready,
	clk,
	reset_n,
	clken,
	phi_inc_i_31,
	phi_inc_i_30,
	phi_inc_i_29,
	phi_inc_i_28,
	phi_inc_i_27,
	phi_inc_i_26,
	phi_inc_i_25,
	phi_inc_i_24,
	phi_inc_i_23,
	phi_inc_i_22,
	phi_inc_i_21,
	phi_inc_i_20,
	phi_inc_i_19,
	phi_inc_i_18,
	phi_inc_i_17,
	phi_inc_i_16,
	phi_inc_i_15,
	phi_inc_i_14,
	phi_inc_i_13,
	phi_inc_i_12,
	phi_inc_i_11,
	phi_inc_i_10,
	phi_inc_i_9,
	phi_inc_i_8,
	phi_inc_i_7,
	phi_inc_i_6,
	phi_inc_i_5,
	phi_inc_i_4,
	phi_inc_i_3,
	phi_inc_i_2,
	phi_inc_i_1,
	phi_inc_i_0)/* synthesis synthesis_greybox=1 */;
output 	sin_o_0;
output 	sin_o_1;
output 	sin_o_2;
output 	sin_o_3;
output 	sin_o_4;
output 	sin_o_5;
output 	sin_o_6;
output 	sin_o_7;
output 	sin_o_8;
output 	sin_o_9;
output 	sin_o_10;
output 	sin_o_11;
output 	sin_o_12;
output 	sin_o_13;
output 	sin_o_14;
output 	sin_o_15;
output 	sin_o_16;
output 	sin_o_17;
output 	cos_o_0;
output 	cos_o_1;
output 	cos_o_2;
output 	cos_o_3;
output 	cos_o_4;
output 	cos_o_5;
output 	cos_o_6;
output 	cos_o_7;
output 	cos_o_8;
output 	cos_o_9;
output 	cos_o_10;
output 	cos_o_11;
output 	cos_o_12;
output 	cos_o_13;
output 	cos_o_14;
output 	cos_o_15;
output 	cos_o_16;
output 	cos_o_17;
output 	data_ready;
input 	clk;
input 	reset_n;
input 	clken;
input 	phi_inc_i_31;
input 	phi_inc_i_30;
input 	phi_inc_i_29;
input 	phi_inc_i_28;
input 	phi_inc_i_27;
input 	phi_inc_i_26;
input 	phi_inc_i_25;
input 	phi_inc_i_24;
input 	phi_inc_i_23;
input 	phi_inc_i_22;
input 	phi_inc_i_21;
input 	phi_inc_i_20;
input 	phi_inc_i_19;
input 	phi_inc_i_18;
input 	phi_inc_i_17;
input 	phi_inc_i_16;
input 	phi_inc_i_15;
input 	phi_inc_i_14;
input 	phi_inc_i_13;
input 	phi_inc_i_12;
input 	phi_inc_i_11;
input 	phi_inc_i_10;
input 	phi_inc_i_9;
input 	phi_inc_i_8;
input 	phi_inc_i_7;
input 	phi_inc_i_6;
input 	phi_inc_i_5;
input 	phi_inc_i_4;
input 	phi_inc_i_3;
input 	phi_inc_i_2;
input 	phi_inc_i_1;
input 	phi_inc_i_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ux005|sin_o[0]~q ;
wire \ux005|sin_o[1]~q ;
wire \ux005|sin_o[2]~q ;
wire \ux005|sin_o[3]~q ;
wire \ux005|sin_o[4]~q ;
wire \ux005|sin_o[5]~q ;
wire \ux005|sin_o[6]~q ;
wire \ux005|sin_o[7]~q ;
wire \ux005|sin_o[8]~q ;
wire \ux005|sin_o[9]~q ;
wire \ux005|sin_o[10]~q ;
wire \ux005|sin_o[11]~q ;
wire \ux005|sin_o[12]~q ;
wire \ux005|sin_o[13]~q ;
wire \ux005|sin_o[14]~q ;
wire \ux005|sin_o[15]~q ;
wire \ux005|sin_o[16]~q ;
wire \ux005|sin_o[17]~q ;
wire \ux005|cos_o[0]~q ;
wire \ux005|cos_o[1]~q ;
wire \ux005|cos_o[2]~q ;
wire \ux005|cos_o[3]~q ;
wire \ux005|cos_o[4]~q ;
wire \ux005|cos_o[5]~q ;
wire \ux005|cos_o[6]~q ;
wire \ux005|cos_o[7]~q ;
wire \ux005|cos_o[8]~q ;
wire \ux005|cos_o[9]~q ;
wire \ux005|cos_o[10]~q ;
wire \ux005|cos_o[11]~q ;
wire \ux005|cos_o[12]~q ;
wire \ux005|cos_o[13]~q ;
wire \ux005|cos_o[14]~q ;
wire \ux005|cos_o[15]~q ;
wire \ux005|cos_o[16]~q ;
wire \ux005|cos_o[17]~q ;
wire \cordinv|cordic_y_res_d[0]~q ;
wire \cordinv|cordic_y_res_2c[0]~q ;
wire \cordinv|cordic_x_res_d[0]~q ;
wire \cordinv|cordic_x_res_2c[0]~q ;
wire \css|seg_rot[1]~q ;
wire \css|seg_rot[0]~q ;
wire \cordinv|cordic_y_res_d[1]~q ;
wire \cordinv|cordic_y_res_2c[1]~q ;
wire \cordinv|cordic_x_res_d[1]~q ;
wire \cordinv|cordic_x_res_2c[1]~q ;
wire \cordinv|cordic_y_res_d[2]~q ;
wire \cordinv|cordic_y_res_2c[2]~q ;
wire \cordinv|cordic_x_res_d[2]~q ;
wire \cordinv|cordic_x_res_2c[2]~q ;
wire \cordinv|cordic_y_res_d[3]~q ;
wire \cordinv|cordic_y_res_2c[3]~q ;
wire \cordinv|cordic_x_res_d[3]~q ;
wire \cordinv|cordic_x_res_2c[3]~q ;
wire \cordinv|cordic_y_res_d[4]~q ;
wire \cordinv|cordic_y_res_2c[4]~q ;
wire \cordinv|cordic_x_res_d[4]~q ;
wire \cordinv|cordic_x_res_2c[4]~q ;
wire \cordinv|cordic_y_res_d[5]~q ;
wire \cordinv|cordic_y_res_2c[5]~q ;
wire \cordinv|cordic_x_res_d[5]~q ;
wire \cordinv|cordic_x_res_2c[5]~q ;
wire \cordinv|cordic_y_res_d[6]~q ;
wire \cordinv|cordic_y_res_2c[6]~q ;
wire \cordinv|cordic_x_res_d[6]~q ;
wire \cordinv|cordic_x_res_2c[6]~q ;
wire \cordinv|cordic_y_res_d[7]~q ;
wire \cordinv|cordic_y_res_2c[7]~q ;
wire \cordinv|cordic_x_res_d[7]~q ;
wire \cordinv|cordic_x_res_2c[7]~q ;
wire \cordinv|cordic_y_res_d[8]~q ;
wire \cordinv|cordic_y_res_2c[8]~q ;
wire \cordinv|cordic_x_res_d[8]~q ;
wire \cordinv|cordic_x_res_2c[8]~q ;
wire \cordinv|cordic_y_res_d[9]~q ;
wire \cordinv|cordic_y_res_2c[9]~q ;
wire \cordinv|cordic_x_res_d[9]~q ;
wire \cordinv|cordic_x_res_2c[9]~q ;
wire \cordinv|cordic_y_res_d[10]~q ;
wire \cordinv|cordic_y_res_2c[10]~q ;
wire \cordinv|cordic_x_res_d[10]~q ;
wire \cordinv|cordic_x_res_2c[10]~q ;
wire \cordinv|cordic_y_res_d[11]~q ;
wire \cordinv|cordic_y_res_2c[11]~q ;
wire \cordinv|cordic_x_res_d[11]~q ;
wire \cordinv|cordic_x_res_2c[11]~q ;
wire \cordinv|cordic_y_res_d[12]~q ;
wire \cordinv|cordic_y_res_2c[12]~q ;
wire \cordinv|cordic_x_res_d[12]~q ;
wire \cordinv|cordic_x_res_2c[12]~q ;
wire \cordinv|cordic_y_res_d[13]~q ;
wire \cordinv|cordic_y_res_2c[13]~q ;
wire \cordinv|cordic_x_res_d[13]~q ;
wire \cordinv|cordic_x_res_2c[13]~q ;
wire \cordinv|cordic_y_res_d[14]~q ;
wire \cordinv|cordic_y_res_2c[14]~q ;
wire \cordinv|cordic_x_res_d[14]~q ;
wire \cordinv|cordic_x_res_2c[14]~q ;
wire \cordinv|cordic_y_res_d[15]~q ;
wire \cordinv|cordic_y_res_2c[15]~q ;
wire \cordinv|cordic_x_res_d[15]~q ;
wire \cordinv|cordic_x_res_2c[15]~q ;
wire \cordinv|cordic_y_res_d[16]~q ;
wire \cordinv|cordic_y_res_2c[16]~q ;
wire \cordinv|cordic_x_res_d[16]~q ;
wire \cordinv|cordic_x_res_2c[16]~q ;
wire \cordinv|cordic_y_res_d[17]~q ;
wire \cordinv|cordic_y_res_2c[17]~q ;
wire \cordinv|cordic_x_res_d[17]~q ;
wire \cordinv|cordic_x_res_2c[17]~q ;
wire \ux002|dxxpdo[20]~q ;
wire \ux002|dxxpdo[19]~q ;
wire \ux001|dxxrv[7]~q ;
wire \u5|a[0]~q ;
wire \u5|xordvalue[11]~q ;
wire \cfs|cor1x[10]~q ;
wire \ux001|dxxrv[6]~q ;
wire \ci|corz[14]~q ;
wire \ux001|dxxrv[5]~q ;
wire \ux002|dxxpdo[18]~q ;
wire \ci|corz[13]~q ;
wire \ux001|dxxrv[4]~q ;
wire \ux002|dxxpdo[17]~q ;
wire \ci|corz[12]~q ;
wire \ux001|dxxrv[3]~q ;
wire \ux002|dxxpdo[16]~q ;
wire \ci|corz[11]~q ;
wire \ux001|dxxrv[2]~q ;
wire \ux002|dxxpdo[15]~q ;
wire \ci|corz[10]~q ;
wire \ux001|dxxrv[1]~q ;
wire \ux002|dxxpdo[14]~q ;
wire \ci|corz[9]~q ;
wire \ux001|dxxrv[0]~q ;
wire \ux002|dxxpdo[13]~q ;
wire \ci|corz[8]~q ;
wire \ux002|dxxpdo[12]~q ;
wire \ci|corz[7]~q ;
wire \ux002|dxxpdo[11]~q ;
wire \ci|corz[6]~q ;
wire \ux002|dxxpdo[10]~q ;
wire \ci|corz[5]~q ;
wire \ux002|dxxpdo[9]~q ;
wire \ci|corz[4]~q ;
wire \ux002|dxxpdo[8]~q ;
wire \ci|corz[3]~q ;
wire \ux002|dxxpdo[7]~q ;
wire \ci|corz[2]~q ;
wire \ux002|dxxpdo[6]~q ;
wire \ci|corz[1]~q ;
wire \ux002|dxxpdo[5]~q ;
wire \ci|corz[0]~q ;
wire \ux002|dxxpdo[4]~q ;
wire \dop|sin_o[0]~0_combout ;
wire \u53|u0|auto_generated|pipeline_dffe[0]~q ;
wire \u52|u0|auto_generated|dffe1~q ;
wire \u53|u0|auto_generated|pipeline_dffe[1]~q ;
wire \u52|u0|auto_generated|dffe2~q ;
wire \u53|u0|auto_generated|pipeline_dffe[2]~q ;
wire \u52|u0|auto_generated|dffe3~q ;
wire \u53|u0|auto_generated|pipeline_dffe[3]~q ;
wire \u52|u0|auto_generated|dffe4~q ;
wire \u53|u0|auto_generated|pipeline_dffe[4]~q ;
wire \u52|u0|auto_generated|dffe5~q ;
wire \u53|u0|auto_generated|pipeline_dffe[5]~q ;
wire \u52|u0|auto_generated|dffe6~q ;
wire \u53|u0|auto_generated|pipeline_dffe[6]~q ;
wire \u52|u0|auto_generated|dffe7~q ;
wire \u53|u0|auto_generated|pipeline_dffe[7]~q ;
wire \u52|u0|auto_generated|dffe8~q ;
wire \u53|u0|auto_generated|pipeline_dffe[8]~q ;
wire \u52|u0|auto_generated|dffe9~q ;
wire \u53|u0|auto_generated|pipeline_dffe[9]~q ;
wire \u52|u0|auto_generated|dffe10~q ;
wire \u53|u0|auto_generated|pipeline_dffe[10]~q ;
wire \u52|u0|auto_generated|dffe11~q ;
wire \u53|u0|auto_generated|pipeline_dffe[11]~q ;
wire \u52|u0|auto_generated|dffe12~q ;
wire \u53|u0|auto_generated|pipeline_dffe[12]~q ;
wire \u52|u0|auto_generated|dffe13~q ;
wire \u53|u0|auto_generated|pipeline_dffe[13]~q ;
wire \u52|u0|auto_generated|dffe14~q ;
wire \u53|u0|auto_generated|pipeline_dffe[14]~q ;
wire \u52|u0|auto_generated|dffe15~q ;
wire \u53|u0|auto_generated|pipeline_dffe[15]~q ;
wire \u52|u0|auto_generated|dffe16~q ;
wire \u53|u0|auto_generated|pipeline_dffe[16]~q ;
wire \u52|u0|auto_generated|dffe17~q ;
wire \u53|u0|auto_generated|pipeline_dffe[17]~q ;
wire \u52|u0|auto_generated|dffe18~q ;
wire \u51|u0|auto_generated|dffe16~q ;
wire \u49|u0|auto_generated|dffe18~q ;
wire \u50|u0|auto_generated|pipeline_dffe[17]~q ;
wire \u50|u0|auto_generated|pipeline_dffe[0]~q ;
wire \u49|u0|auto_generated|dffe1~q ;
wire \u50|u0|auto_generated|pipeline_dffe[1]~q ;
wire \u49|u0|auto_generated|dffe2~q ;
wire \u50|u0|auto_generated|pipeline_dffe[2]~q ;
wire \u49|u0|auto_generated|dffe3~q ;
wire \u50|u0|auto_generated|pipeline_dffe[3]~q ;
wire \u49|u0|auto_generated|dffe4~q ;
wire \u50|u0|auto_generated|pipeline_dffe[4]~q ;
wire \u49|u0|auto_generated|dffe5~q ;
wire \u50|u0|auto_generated|pipeline_dffe[5]~q ;
wire \u49|u0|auto_generated|dffe6~q ;
wire \u50|u0|auto_generated|pipeline_dffe[6]~q ;
wire \u49|u0|auto_generated|dffe7~q ;
wire \u50|u0|auto_generated|pipeline_dffe[7]~q ;
wire \u49|u0|auto_generated|dffe8~q ;
wire \u50|u0|auto_generated|pipeline_dffe[8]~q ;
wire \u49|u0|auto_generated|dffe9~q ;
wire \u50|u0|auto_generated|pipeline_dffe[9]~q ;
wire \u49|u0|auto_generated|dffe10~q ;
wire \u50|u0|auto_generated|pipeline_dffe[10]~q ;
wire \u49|u0|auto_generated|dffe11~q ;
wire \u50|u0|auto_generated|pipeline_dffe[11]~q ;
wire \u49|u0|auto_generated|dffe12~q ;
wire \u50|u0|auto_generated|pipeline_dffe[12]~q ;
wire \u49|u0|auto_generated|dffe13~q ;
wire \u50|u0|auto_generated|pipeline_dffe[13]~q ;
wire \u49|u0|auto_generated|dffe14~q ;
wire \u50|u0|auto_generated|pipeline_dffe[14]~q ;
wire \u49|u0|auto_generated|dffe15~q ;
wire \u50|u0|auto_generated|pipeline_dffe[15]~q ;
wire \u49|u0|auto_generated|dffe16~q ;
wire \u50|u0|auto_generated|pipeline_dffe[16]~q ;
wire \u49|u0|auto_generated|dffe17~q ;
wire \u48|u0|auto_generated|dffe16~q ;
wire \u47|u0|auto_generated|pipeline_dffe[17]~q ;
wire \u46|u0|auto_generated|dffe18~q ;
wire \u46|u0|auto_generated|dffe17~q ;
wire \u47|u0|auto_generated|pipeline_dffe[16]~q ;
wire \u47|u0|auto_generated|pipeline_dffe[0]~q ;
wire \u48|u0|auto_generated|dffe15~q ;
wire \u46|u0|auto_generated|dffe1~q ;
wire \u47|u0|auto_generated|pipeline_dffe[1]~q ;
wire \u46|u0|auto_generated|dffe2~q ;
wire \u47|u0|auto_generated|pipeline_dffe[2]~q ;
wire \u46|u0|auto_generated|dffe3~q ;
wire \u47|u0|auto_generated|pipeline_dffe[3]~q ;
wire \u46|u0|auto_generated|dffe4~q ;
wire \u47|u0|auto_generated|pipeline_dffe[4]~q ;
wire \u46|u0|auto_generated|dffe5~q ;
wire \u47|u0|auto_generated|pipeline_dffe[5]~q ;
wire \u46|u0|auto_generated|dffe6~q ;
wire \u47|u0|auto_generated|pipeline_dffe[6]~q ;
wire \u46|u0|auto_generated|dffe7~q ;
wire \u47|u0|auto_generated|pipeline_dffe[7]~q ;
wire \u46|u0|auto_generated|dffe8~q ;
wire \u47|u0|auto_generated|pipeline_dffe[8]~q ;
wire \u46|u0|auto_generated|dffe9~q ;
wire \u47|u0|auto_generated|pipeline_dffe[9]~q ;
wire \u46|u0|auto_generated|dffe10~q ;
wire \u47|u0|auto_generated|pipeline_dffe[10]~q ;
wire \u46|u0|auto_generated|dffe11~q ;
wire \u47|u0|auto_generated|pipeline_dffe[11]~q ;
wire \u46|u0|auto_generated|dffe12~q ;
wire \u47|u0|auto_generated|pipeline_dffe[12]~q ;
wire \u46|u0|auto_generated|dffe13~q ;
wire \u47|u0|auto_generated|pipeline_dffe[13]~q ;
wire \u46|u0|auto_generated|dffe14~q ;
wire \u47|u0|auto_generated|pipeline_dffe[14]~q ;
wire \u46|u0|auto_generated|dffe15~q ;
wire \u47|u0|auto_generated|pipeline_dffe[15]~q ;
wire \u46|u0|auto_generated|dffe16~q ;
wire \u48|u0|auto_generated|dffe14~q ;
wire \u45|u0|auto_generated|dffe16~q ;
wire \u43|u0|auto_generated|dffe18~q ;
wire \u44|u0|auto_generated|pipeline_dffe[17]~q ;
wire \u48|u0|auto_generated|dffe13~q ;
wire \u43|u0|auto_generated|dffe16~q ;
wire \u43|u0|auto_generated|dffe17~q ;
wire \u48|u0|auto_generated|dffe12~q ;
wire \u45|u0|auto_generated|dffe15~q ;
wire \u44|u0|auto_generated|pipeline_dffe[16]~q ;
wire \u44|u0|auto_generated|pipeline_dffe[15]~q ;
wire \u44|u0|auto_generated|pipeline_dffe[0]~q ;
wire \u48|u0|auto_generated|dffe11~q ;
wire \u45|u0|auto_generated|dffe14~q ;
wire \u42|u0|auto_generated|dffe16~q ;
wire \u41|u0|auto_generated|pipeline_dffe[17]~q ;
wire \u43|u0|auto_generated|dffe1~q ;
wire \u40|u0|auto_generated|dffe18~q ;
wire \u44|u0|auto_generated|pipeline_dffe[1]~q ;
wire \u43|u0|auto_generated|dffe2~q ;
wire \u44|u0|auto_generated|pipeline_dffe[2]~q ;
wire \u43|u0|auto_generated|dffe3~q ;
wire \u44|u0|auto_generated|pipeline_dffe[3]~q ;
wire \u43|u0|auto_generated|dffe4~q ;
wire \u44|u0|auto_generated|pipeline_dffe[4]~q ;
wire \u43|u0|auto_generated|dffe5~q ;
wire \u44|u0|auto_generated|pipeline_dffe[5]~q ;
wire \u43|u0|auto_generated|dffe6~q ;
wire \u44|u0|auto_generated|pipeline_dffe[6]~q ;
wire \u43|u0|auto_generated|dffe7~q ;
wire \u44|u0|auto_generated|pipeline_dffe[7]~q ;
wire \u43|u0|auto_generated|dffe8~q ;
wire \u44|u0|auto_generated|pipeline_dffe[8]~q ;
wire \u43|u0|auto_generated|dffe9~q ;
wire \u44|u0|auto_generated|pipeline_dffe[9]~q ;
wire \u43|u0|auto_generated|dffe10~q ;
wire \u44|u0|auto_generated|pipeline_dffe[10]~q ;
wire \u43|u0|auto_generated|dffe11~q ;
wire \u44|u0|auto_generated|pipeline_dffe[11]~q ;
wire \u43|u0|auto_generated|dffe12~q ;
wire \u44|u0|auto_generated|pipeline_dffe[12]~q ;
wire \u43|u0|auto_generated|dffe13~q ;
wire \u44|u0|auto_generated|pipeline_dffe[13]~q ;
wire \u43|u0|auto_generated|dffe14~q ;
wire \u44|u0|auto_generated|pipeline_dffe[14]~q ;
wire \u43|u0|auto_generated|dffe15~q ;
wire \u48|u0|auto_generated|dffe10~q ;
wire \u45|u0|auto_generated|dffe13~q ;
wire \u48|u0|auto_generated|dffe9~q ;
wire \u45|u0|auto_generated|dffe12~q ;
wire \u42|u0|auto_generated|dffe15~q ;
wire \u40|u0|auto_generated|dffe17~q ;
wire \u41|u0|auto_generated|pipeline_dffe[16]~q ;
wire \u40|u0|auto_generated|dffe15~q ;
wire \u40|u0|auto_generated|dffe16~q ;
wire \u48|u0|auto_generated|dffe8~q ;
wire \u45|u0|auto_generated|dffe11~q ;
wire \u42|u0|auto_generated|dffe14~q ;
wire \u39|u0|auto_generated|dffe16~q ;
wire \u37|u0|auto_generated|dffe18~q ;
wire \u41|u0|auto_generated|pipeline_dffe[14]~q ;
wire \u41|u0|auto_generated|pipeline_dffe[15]~q ;
wire \u38|u0|auto_generated|pipeline_dffe[17]~q ;
wire \u41|u0|auto_generated|pipeline_dffe[0]~q ;
wire \u48|u0|auto_generated|dffe7~q ;
wire \u45|u0|auto_generated|dffe10~q ;
wire \u42|u0|auto_generated|dffe13~q ;
wire \u40|u0|auto_generated|dffe1~q ;
wire \u41|u0|auto_generated|pipeline_dffe[1]~q ;
wire \u40|u0|auto_generated|dffe2~q ;
wire \u41|u0|auto_generated|pipeline_dffe[2]~q ;
wire \u40|u0|auto_generated|dffe3~q ;
wire \u41|u0|auto_generated|pipeline_dffe[3]~q ;
wire \u40|u0|auto_generated|dffe4~q ;
wire \u41|u0|auto_generated|pipeline_dffe[4]~q ;
wire \u40|u0|auto_generated|dffe5~q ;
wire \u41|u0|auto_generated|pipeline_dffe[5]~q ;
wire \u40|u0|auto_generated|dffe6~q ;
wire \u41|u0|auto_generated|pipeline_dffe[6]~q ;
wire \u40|u0|auto_generated|dffe7~q ;
wire \u41|u0|auto_generated|pipeline_dffe[7]~q ;
wire \u40|u0|auto_generated|dffe8~q ;
wire \u41|u0|auto_generated|pipeline_dffe[8]~q ;
wire \u40|u0|auto_generated|dffe9~q ;
wire \u41|u0|auto_generated|pipeline_dffe[9]~q ;
wire \u40|u0|auto_generated|dffe10~q ;
wire \u41|u0|auto_generated|pipeline_dffe[10]~q ;
wire \u40|u0|auto_generated|dffe11~q ;
wire \u41|u0|auto_generated|pipeline_dffe[11]~q ;
wire \u40|u0|auto_generated|dffe12~q ;
wire \u41|u0|auto_generated|pipeline_dffe[12]~q ;
wire \u40|u0|auto_generated|dffe13~q ;
wire \u41|u0|auto_generated|pipeline_dffe[13]~q ;
wire \u40|u0|auto_generated|dffe14~q ;
wire \u48|u0|auto_generated|dffe6~q ;
wire \u45|u0|auto_generated|dffe9~q ;
wire \u42|u0|auto_generated|dffe12~q ;
wire \u39|u0|auto_generated|dffe15~q ;
wire \u38|u0|auto_generated|pipeline_dffe[16]~q ;
wire \u37|u0|auto_generated|dffe17~q ;
wire \u48|u0|auto_generated|dffe5~q ;
wire \u45|u0|auto_generated|dffe8~q ;
wire \u42|u0|auto_generated|dffe11~q ;
wire \u39|u0|auto_generated|dffe14~q ;
wire \u36|u0|auto_generated|dffe16~q ;
wire \u38|u0|auto_generated|pipeline_dffe[15]~q ;
wire \u35|u0|auto_generated|pipeline_dffe[17]~q ;
wire \u37|u0|auto_generated|dffe16~q ;
wire \u34|u0|auto_generated|dffe18~q ;
wire \u37|u0|auto_generated|dffe14~q ;
wire \u37|u0|auto_generated|dffe15~q ;
wire \u48|u0|auto_generated|dffe4~q ;
wire \u45|u0|auto_generated|dffe7~q ;
wire \u42|u0|auto_generated|dffe10~q ;
wire \u39|u0|auto_generated|dffe13~q ;
wire \u38|u0|auto_generated|pipeline_dffe[14]~q ;
wire \u38|u0|auto_generated|pipeline_dffe[13]~q ;
wire \u38|u0|auto_generated|pipeline_dffe[0]~q ;
wire \u48|u0|auto_generated|dffe3~q ;
wire \u45|u0|auto_generated|dffe6~q ;
wire \u42|u0|auto_generated|dffe9~q ;
wire \u39|u0|auto_generated|dffe12~q ;
wire \u36|u0|auto_generated|dffe15~q ;
wire \u34|u0|auto_generated|dffe17~q ;
wire \u37|u0|auto_generated|dffe1~q ;
wire \u35|u0|auto_generated|pipeline_dffe[16]~q ;
wire \u38|u0|auto_generated|pipeline_dffe[1]~q ;
wire \u37|u0|auto_generated|dffe2~q ;
wire \u38|u0|auto_generated|pipeline_dffe[2]~q ;
wire \u37|u0|auto_generated|dffe3~q ;
wire \u38|u0|auto_generated|pipeline_dffe[3]~q ;
wire \u37|u0|auto_generated|dffe4~q ;
wire \u38|u0|auto_generated|pipeline_dffe[4]~q ;
wire \u37|u0|auto_generated|dffe5~q ;
wire \u38|u0|auto_generated|pipeline_dffe[5]~q ;
wire \u37|u0|auto_generated|dffe6~q ;
wire \u38|u0|auto_generated|pipeline_dffe[6]~q ;
wire \u37|u0|auto_generated|dffe7~q ;
wire \u38|u0|auto_generated|pipeline_dffe[7]~q ;
wire \u37|u0|auto_generated|dffe8~q ;
wire \u38|u0|auto_generated|pipeline_dffe[8]~q ;
wire \u37|u0|auto_generated|dffe9~q ;
wire \u38|u0|auto_generated|pipeline_dffe[9]~q ;
wire \u37|u0|auto_generated|dffe10~q ;
wire \u38|u0|auto_generated|pipeline_dffe[10]~q ;
wire \u37|u0|auto_generated|dffe11~q ;
wire \u38|u0|auto_generated|pipeline_dffe[11]~q ;
wire \u37|u0|auto_generated|dffe12~q ;
wire \u38|u0|auto_generated|pipeline_dffe[12]~q ;
wire \u37|u0|auto_generated|dffe13~q ;
wire \u48|u0|auto_generated|dffe2~q ;
wire \u45|u0|auto_generated|dffe5~q ;
wire \u42|u0|auto_generated|dffe8~q ;
wire \u39|u0|auto_generated|dffe11~q ;
wire \u36|u0|auto_generated|dffe14~q ;
wire \u33|u0|auto_generated|dffe16~q ;
wire \u34|u0|auto_generated|dffe16~q ;
wire \u31|u0|auto_generated|dffe18~q ;
wire \u35|u0|auto_generated|pipeline_dffe[15]~q ;
wire \u32|u0|auto_generated|pipeline_dffe[17]~q ;
wire \u48|u0|auto_generated|dffe1~q ;
wire \u45|u0|auto_generated|dffe4~q ;
wire \u42|u0|auto_generated|dffe7~q ;
wire \u39|u0|auto_generated|dffe10~q ;
wire \u36|u0|auto_generated|dffe13~q ;
wire \u34|u0|auto_generated|dffe15~q ;
wire \u35|u0|auto_generated|pipeline_dffe[14]~q ;
wire \u34|u0|auto_generated|dffe13~q ;
wire \u34|u0|auto_generated|dffe14~q ;
wire \u45|u0|auto_generated|dffe3~q ;
wire \u42|u0|auto_generated|dffe6~q ;
wire \u39|u0|auto_generated|dffe9~q ;
wire \u36|u0|auto_generated|dffe12~q ;
wire \u33|u0|auto_generated|dffe15~q ;
wire \u32|u0|auto_generated|pipeline_dffe[16]~q ;
wire \u35|u0|auto_generated|pipeline_dffe[12]~q ;
wire \u35|u0|auto_generated|pipeline_dffe[13]~q ;
wire \u31|u0|auto_generated|dffe17~q ;
wire \u35|u0|auto_generated|pipeline_dffe[0]~q ;
wire \u45|u0|auto_generated|dffe2~q ;
wire \u42|u0|auto_generated|dffe5~q ;
wire \u39|u0|auto_generated|dffe8~q ;
wire \u36|u0|auto_generated|dffe11~q ;
wire \u33|u0|auto_generated|dffe14~q ;
wire \u30|u0|auto_generated|dffe16~q ;
wire \u32|u0|auto_generated|pipeline_dffe[15]~q ;
wire \u29|u0|auto_generated|pipeline_dffe[17]~q ;
wire \u34|u0|auto_generated|dffe1~q ;
wire \u31|u0|auto_generated|dffe16~q ;
wire \u28|u0|auto_generated|dffe18~q ;
wire \u35|u0|auto_generated|pipeline_dffe[1]~q ;
wire \u34|u0|auto_generated|dffe2~q ;
wire \u35|u0|auto_generated|pipeline_dffe[2]~q ;
wire \u34|u0|auto_generated|dffe3~q ;
wire \u35|u0|auto_generated|pipeline_dffe[3]~q ;
wire \u34|u0|auto_generated|dffe4~q ;
wire \u35|u0|auto_generated|pipeline_dffe[4]~q ;
wire \u34|u0|auto_generated|dffe5~q ;
wire \u35|u0|auto_generated|pipeline_dffe[5]~q ;
wire \u34|u0|auto_generated|dffe6~q ;
wire \u35|u0|auto_generated|pipeline_dffe[6]~q ;
wire \u34|u0|auto_generated|dffe7~q ;
wire \u35|u0|auto_generated|pipeline_dffe[7]~q ;
wire \u34|u0|auto_generated|dffe8~q ;
wire \u35|u0|auto_generated|pipeline_dffe[8]~q ;
wire \u34|u0|auto_generated|dffe9~q ;
wire \u35|u0|auto_generated|pipeline_dffe[9]~q ;
wire \u34|u0|auto_generated|dffe10~q ;
wire \u35|u0|auto_generated|pipeline_dffe[10]~q ;
wire \u34|u0|auto_generated|dffe11~q ;
wire \u35|u0|auto_generated|pipeline_dffe[11]~q ;
wire \u34|u0|auto_generated|dffe12~q ;
wire \u45|u0|auto_generated|dffe1~q ;
wire \u42|u0|auto_generated|dffe4~q ;
wire \u39|u0|auto_generated|dffe7~q ;
wire \u36|u0|auto_generated|dffe10~q ;
wire \u33|u0|auto_generated|dffe13~q ;
wire \u32|u0|auto_generated|pipeline_dffe[14]~q ;
wire \u31|u0|auto_generated|dffe15~q ;
wire \u42|u0|auto_generated|dffe3~q ;
wire \u39|u0|auto_generated|dffe6~q ;
wire \u36|u0|auto_generated|dffe9~q ;
wire \u33|u0|auto_generated|dffe12~q ;
wire \u30|u0|auto_generated|dffe15~q ;
wire \u32|u0|auto_generated|pipeline_dffe[13]~q ;
wire \u28|u0|auto_generated|dffe17~q ;
wire \u31|u0|auto_generated|dffe14~q ;
wire \u29|u0|auto_generated|pipeline_dffe[16]~q ;
wire \u31|u0|auto_generated|dffe12~q ;
wire \u31|u0|auto_generated|dffe13~q ;
wire \u42|u0|auto_generated|dffe2~q ;
wire \u39|u0|auto_generated|dffe5~q ;
wire \u36|u0|auto_generated|dffe8~q ;
wire \u33|u0|auto_generated|dffe11~q ;
wire \u30|u0|auto_generated|dffe14~q ;
wire \u27|u0|auto_generated|dffe16~q ;
wire \u32|u0|auto_generated|pipeline_dffe[12]~q ;
wire \u28|u0|auto_generated|dffe16~q ;
wire \u25|u0|auto_generated|dffe18~q ;
wire \u32|u0|auto_generated|pipeline_dffe[11]~q ;
wire \u29|u0|auto_generated|pipeline_dffe[15]~q ;
wire \u26|u0|auto_generated|pipeline_dffe[17]~q ;
wire \u32|u0|auto_generated|pipeline_dffe[0]~q ;
wire \u42|u0|auto_generated|dffe1~q ;
wire \u39|u0|auto_generated|dffe4~q ;
wire \u36|u0|auto_generated|dffe7~q ;
wire \u33|u0|auto_generated|dffe10~q ;
wire \u30|u0|auto_generated|dffe13~q ;
wire \u28|u0|auto_generated|dffe15~q ;
wire \u31|u0|auto_generated|dffe1~q ;
wire \u29|u0|auto_generated|pipeline_dffe[14]~q ;
wire \u32|u0|auto_generated|pipeline_dffe[1]~q ;
wire \u31|u0|auto_generated|dffe2~q ;
wire \u32|u0|auto_generated|pipeline_dffe[2]~q ;
wire \u31|u0|auto_generated|dffe3~q ;
wire \u32|u0|auto_generated|pipeline_dffe[3]~q ;
wire \u31|u0|auto_generated|dffe4~q ;
wire \u32|u0|auto_generated|pipeline_dffe[4]~q ;
wire \u31|u0|auto_generated|dffe5~q ;
wire \u32|u0|auto_generated|pipeline_dffe[5]~q ;
wire \u31|u0|auto_generated|dffe6~q ;
wire \u32|u0|auto_generated|pipeline_dffe[6]~q ;
wire \u31|u0|auto_generated|dffe7~q ;
wire \u32|u0|auto_generated|pipeline_dffe[7]~q ;
wire \u31|u0|auto_generated|dffe8~q ;
wire \u32|u0|auto_generated|pipeline_dffe[8]~q ;
wire \u31|u0|auto_generated|dffe9~q ;
wire \u32|u0|auto_generated|pipeline_dffe[9]~q ;
wire \u31|u0|auto_generated|dffe10~q ;
wire \u32|u0|auto_generated|pipeline_dffe[10]~q ;
wire \u31|u0|auto_generated|dffe11~q ;
wire \u39|u0|auto_generated|dffe3~q ;
wire \u36|u0|auto_generated|dffe6~q ;
wire \u33|u0|auto_generated|dffe9~q ;
wire \u30|u0|auto_generated|dffe12~q ;
wire \u27|u0|auto_generated|dffe15~q ;
wire \u28|u0|auto_generated|dffe14~q ;
wire \u26|u0|auto_generated|pipeline_dffe[16]~q ;
wire \u29|u0|auto_generated|pipeline_dffe[13]~q ;
wire \u25|u0|auto_generated|dffe17~q ;
wire \u39|u0|auto_generated|dffe2~q ;
wire \u36|u0|auto_generated|dffe5~q ;
wire \u33|u0|auto_generated|dffe8~q ;
wire \u30|u0|auto_generated|dffe11~q ;
wire \u27|u0|auto_generated|dffe14~q ;
wire \u24|u0|auto_generated|dffe16~q ;
wire \u28|u0|auto_generated|dffe13~q ;
wire \u26|u0|auto_generated|pipeline_dffe[15]~q ;
wire \u23|u0|auto_generated|pipeline_dffe[17]~q ;
wire \u29|u0|auto_generated|pipeline_dffe[12]~q ;
wire \u25|u0|auto_generated|dffe16~q ;
wire \u22|u0|auto_generated|dffe18~q ;
wire \u28|u0|auto_generated|dffe11~q ;
wire \u28|u0|auto_generated|dffe12~q ;
wire \u39|u0|auto_generated|dffe1~q ;
wire \u36|u0|auto_generated|dffe4~q ;
wire \u33|u0|auto_generated|dffe7~q ;
wire \u30|u0|auto_generated|dffe10~q ;
wire \u27|u0|auto_generated|dffe13~q ;
wire \u26|u0|auto_generated|pipeline_dffe[14]~q ;
wire \u29|u0|auto_generated|pipeline_dffe[10]~q ;
wire \u29|u0|auto_generated|pipeline_dffe[11]~q ;
wire \u25|u0|auto_generated|dffe15~q ;
wire \u29|u0|auto_generated|pipeline_dffe[0]~q ;
wire \u36|u0|auto_generated|dffe3~q ;
wire \u33|u0|auto_generated|dffe6~q ;
wire \u30|u0|auto_generated|dffe9~q ;
wire \u27|u0|auto_generated|dffe12~q ;
wire \u24|u0|auto_generated|dffe15~q ;
wire \u26|u0|auto_generated|pipeline_dffe[13]~q ;
wire \u22|u0|auto_generated|dffe17~q ;
wire \u28|u0|auto_generated|dffe1~q ;
wire \u25|u0|auto_generated|dffe14~q ;
wire \u23|u0|auto_generated|pipeline_dffe[16]~q ;
wire \u29|u0|auto_generated|pipeline_dffe[1]~q ;
wire \u28|u0|auto_generated|dffe2~q ;
wire \u29|u0|auto_generated|pipeline_dffe[2]~q ;
wire \u28|u0|auto_generated|dffe3~q ;
wire \u29|u0|auto_generated|pipeline_dffe[3]~q ;
wire \u28|u0|auto_generated|dffe4~q ;
wire \u29|u0|auto_generated|pipeline_dffe[4]~q ;
wire \u28|u0|auto_generated|dffe5~q ;
wire \u29|u0|auto_generated|pipeline_dffe[5]~q ;
wire \u28|u0|auto_generated|dffe6~q ;
wire \u29|u0|auto_generated|pipeline_dffe[6]~q ;
wire \u28|u0|auto_generated|dffe7~q ;
wire \u29|u0|auto_generated|pipeline_dffe[7]~q ;
wire \u28|u0|auto_generated|dffe8~q ;
wire \u29|u0|auto_generated|pipeline_dffe[8]~q ;
wire \u28|u0|auto_generated|dffe9~q ;
wire \u29|u0|auto_generated|pipeline_dffe[9]~q ;
wire \u28|u0|auto_generated|dffe10~q ;
wire \u36|u0|auto_generated|dffe2~q ;
wire \u33|u0|auto_generated|dffe5~q ;
wire \u30|u0|auto_generated|dffe8~q ;
wire \u27|u0|auto_generated|dffe11~q ;
wire \u24|u0|auto_generated|dffe14~q ;
wire \u21|u0|auto_generated|dffe16~q ;
wire \u26|u0|auto_generated|pipeline_dffe[12]~q ;
wire \u22|u0|auto_generated|dffe16~q ;
wire \u19|u0|auto_generated|dffe18~q ;
wire \u25|u0|auto_generated|dffe13~q ;
wire \u23|u0|auto_generated|pipeline_dffe[15]~q ;
wire \u20|u0|auto_generated|pipeline_dffe[17]~q ;
wire \u36|u0|auto_generated|dffe1~q ;
wire \u33|u0|auto_generated|dffe4~q ;
wire \u30|u0|auto_generated|dffe7~q ;
wire \u27|u0|auto_generated|dffe10~q ;
wire \u24|u0|auto_generated|dffe13~q ;
wire \u26|u0|auto_generated|pipeline_dffe[11]~q ;
wire \u22|u0|auto_generated|dffe15~q ;
wire \u25|u0|auto_generated|dffe12~q ;
wire \u23|u0|auto_generated|pipeline_dffe[14]~q ;
wire \u25|u0|auto_generated|dffe10~q ;
wire \u25|u0|auto_generated|dffe11~q ;
wire \u33|u0|auto_generated|dffe3~q ;
wire \u30|u0|auto_generated|dffe6~q ;
wire \u27|u0|auto_generated|dffe9~q ;
wire \u24|u0|auto_generated|dffe12~q ;
wire \u21|u0|auto_generated|dffe15~q ;
wire \u26|u0|auto_generated|pipeline_dffe[10]~q ;
wire \u22|u0|auto_generated|dffe14~q ;
wire \u20|u0|auto_generated|pipeline_dffe[16]~q ;
wire \u26|u0|auto_generated|pipeline_dffe[9]~q ;
wire \u23|u0|auto_generated|pipeline_dffe[13]~q ;
wire \u19|u0|auto_generated|dffe17~q ;
wire \u26|u0|auto_generated|pipeline_dffe[0]~q ;
wire \u33|u0|auto_generated|dffe2~q ;
wire \u30|u0|auto_generated|dffe5~q ;
wire \u27|u0|auto_generated|dffe8~q ;
wire \u24|u0|auto_generated|dffe11~q ;
wire \u21|u0|auto_generated|dffe14~q ;
wire \u18|u0|auto_generated|dffe16~q ;
wire \u22|u0|auto_generated|dffe13~q ;
wire \u20|u0|auto_generated|pipeline_dffe[15]~q ;
wire \u17|u0|auto_generated|pipeline_dffe[17]~q ;
wire \u25|u0|auto_generated|dffe1~q ;
wire \u23|u0|auto_generated|pipeline_dffe[12]~q ;
wire \u19|u0|auto_generated|dffe16~q ;
wire \u16|u0|auto_generated|dffe18~q ;
wire \u26|u0|auto_generated|pipeline_dffe[1]~q ;
wire \u25|u0|auto_generated|dffe2~q ;
wire \u26|u0|auto_generated|pipeline_dffe[2]~q ;
wire \u25|u0|auto_generated|dffe3~q ;
wire \u26|u0|auto_generated|pipeline_dffe[3]~q ;
wire \u25|u0|auto_generated|dffe4~q ;
wire \u26|u0|auto_generated|pipeline_dffe[4]~q ;
wire \u25|u0|auto_generated|dffe5~q ;
wire \u26|u0|auto_generated|pipeline_dffe[5]~q ;
wire \u25|u0|auto_generated|dffe6~q ;
wire \u26|u0|auto_generated|pipeline_dffe[6]~q ;
wire \u25|u0|auto_generated|dffe7~q ;
wire \u26|u0|auto_generated|pipeline_dffe[7]~q ;
wire \u25|u0|auto_generated|dffe8~q ;
wire \u26|u0|auto_generated|pipeline_dffe[8]~q ;
wire \u25|u0|auto_generated|dffe9~q ;
wire \u33|u0|auto_generated|dffe1~q ;
wire \u30|u0|auto_generated|dffe4~q ;
wire \u27|u0|auto_generated|dffe7~q ;
wire \u24|u0|auto_generated|dffe10~q ;
wire \u21|u0|auto_generated|dffe13~q ;
wire \u22|u0|auto_generated|dffe12~q ;
wire \u20|u0|auto_generated|pipeline_dffe[14]~q ;
wire \u23|u0|auto_generated|pipeline_dffe[11]~q ;
wire \u19|u0|auto_generated|dffe15~q ;
wire \u30|u0|auto_generated|dffe3~q ;
wire \u27|u0|auto_generated|dffe6~q ;
wire \u24|u0|auto_generated|dffe9~q ;
wire \u21|u0|auto_generated|dffe12~q ;
wire \u18|u0|auto_generated|dffe15~q ;
wire \u22|u0|auto_generated|dffe11~q ;
wire \u20|u0|auto_generated|pipeline_dffe[13]~q ;
wire \u16|u0|auto_generated|dffe17~q ;
wire \u23|u0|auto_generated|pipeline_dffe[10]~q ;
wire \u19|u0|auto_generated|dffe14~q ;
wire \u17|u0|auto_generated|pipeline_dffe[16]~q ;
wire \u22|u0|auto_generated|dffe9~q ;
wire \u22|u0|auto_generated|dffe10~q ;
wire \u30|u0|auto_generated|dffe2~q ;
wire \u27|u0|auto_generated|dffe5~q ;
wire \u24|u0|auto_generated|dffe8~q ;
wire \u21|u0|auto_generated|dffe11~q ;
wire \u18|u0|auto_generated|dffe14~q ;
wire \u15|u0|auto_generated|dffe16~q ;
wire \u20|u0|auto_generated|pipeline_dffe[12]~q ;
wire \u16|u0|auto_generated|dffe16~q ;
wire \u13|u0|auto_generated|dffe18~q ;
wire \u23|u0|auto_generated|pipeline_dffe[8]~q ;
wire \u23|u0|auto_generated|pipeline_dffe[9]~q ;
wire \u19|u0|auto_generated|dffe13~q ;
wire \u17|u0|auto_generated|pipeline_dffe[15]~q ;
wire \u14|u0|auto_generated|pipeline_dffe[17]~q ;
wire \u23|u0|auto_generated|pipeline_dffe[0]~q ;
wire \u30|u0|auto_generated|dffe1~q ;
wire \u27|u0|auto_generated|dffe4~q ;
wire \u24|u0|auto_generated|dffe7~q ;
wire \u21|u0|auto_generated|dffe10~q ;
wire \u18|u0|auto_generated|dffe13~q ;
wire \u20|u0|auto_generated|pipeline_dffe[11]~q ;
wire \u16|u0|auto_generated|dffe15~q ;
wire \u22|u0|auto_generated|dffe1~q ;
wire \u19|u0|auto_generated|dffe12~q ;
wire \u17|u0|auto_generated|pipeline_dffe[14]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[31]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[30]~q ;
wire \u23|u0|auto_generated|pipeline_dffe[1]~q ;
wire \u22|u0|auto_generated|dffe2~q ;
wire \u23|u0|auto_generated|pipeline_dffe[2]~q ;
wire \u22|u0|auto_generated|dffe3~q ;
wire \u23|u0|auto_generated|pipeline_dffe[3]~q ;
wire \u22|u0|auto_generated|dffe4~q ;
wire \u23|u0|auto_generated|pipeline_dffe[4]~q ;
wire \u22|u0|auto_generated|dffe5~q ;
wire \u23|u0|auto_generated|pipeline_dffe[5]~q ;
wire \u22|u0|auto_generated|dffe6~q ;
wire \u23|u0|auto_generated|pipeline_dffe[6]~q ;
wire \u22|u0|auto_generated|dffe7~q ;
wire \u23|u0|auto_generated|pipeline_dffe[7]~q ;
wire \u22|u0|auto_generated|dffe8~q ;
wire \u27|u0|auto_generated|dffe3~q ;
wire \u24|u0|auto_generated|dffe6~q ;
wire \u21|u0|auto_generated|dffe9~q ;
wire \u18|u0|auto_generated|dffe12~q ;
wire \u15|u0|auto_generated|dffe15~q ;
wire \u20|u0|auto_generated|pipeline_dffe[10]~q ;
wire \u16|u0|auto_generated|dffe14~q ;
wire \u14|u0|auto_generated|pipeline_dffe[16]~q ;
wire \u19|u0|auto_generated|dffe11~q ;
wire \u17|u0|auto_generated|pipeline_dffe[13]~q ;
wire \u13|u0|auto_generated|dffe17~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[29]~q ;
wire \u27|u0|auto_generated|dffe2~q ;
wire \u24|u0|auto_generated|dffe5~q ;
wire \u21|u0|auto_generated|dffe8~q ;
wire \u18|u0|auto_generated|dffe11~q ;
wire \u15|u0|auto_generated|dffe14~q ;
wire \u12|u0|auto_generated|dffe16~q ;
wire \u20|u0|auto_generated|pipeline_dffe[9]~q ;
wire \u16|u0|auto_generated|dffe13~q ;
wire \u14|u0|auto_generated|pipeline_dffe[15]~q ;
wire \u11|u0|auto_generated|pipeline_dffe[17]~q ;
wire \u19|u0|auto_generated|dffe10~q ;
wire \u17|u0|auto_generated|pipeline_dffe[12]~q ;
wire \u13|u0|auto_generated|dffe16~q ;
wire \u10|u0|auto_generated|dffe18~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[28]~q ;
wire \u19|u0|auto_generated|dffe8~q ;
wire \u19|u0|auto_generated|dffe9~q ;
wire \u27|u0|auto_generated|dffe1~q ;
wire \u24|u0|auto_generated|dffe4~q ;
wire \u21|u0|auto_generated|dffe7~q ;
wire \u18|u0|auto_generated|dffe10~q ;
wire \u15|u0|auto_generated|dffe13~q ;
wire \u20|u0|auto_generated|pipeline_dffe[8]~q ;
wire \u16|u0|auto_generated|dffe12~q ;
wire \u14|u0|auto_generated|pipeline_dffe[14]~q ;
wire \u20|u0|auto_generated|pipeline_dffe[7]~q ;
wire \u17|u0|auto_generated|pipeline_dffe[11]~q ;
wire \u13|u0|auto_generated|dffe15~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[27]~q ;
wire \u20|u0|auto_generated|pipeline_dffe[0]~q ;
wire \u24|u0|auto_generated|dffe3~q ;
wire \u21|u0|auto_generated|dffe6~q ;
wire \u18|u0|auto_generated|dffe9~q ;
wire \u15|u0|auto_generated|dffe12~q ;
wire \u12|u0|auto_generated|dffe15~q ;
wire \u16|u0|auto_generated|dffe11~q ;
wire \u14|u0|auto_generated|pipeline_dffe[13]~q ;
wire \u10|u0|auto_generated|dffe17~q ;
wire \u19|u0|auto_generated|dffe1~q ;
wire \u17|u0|auto_generated|pipeline_dffe[10]~q ;
wire \u13|u0|auto_generated|dffe14~q ;
wire \u11|u0|auto_generated|pipeline_dffe[16]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[26]~q ;
wire \u20|u0|auto_generated|pipeline_dffe[1]~q ;
wire \u19|u0|auto_generated|dffe2~q ;
wire \u20|u0|auto_generated|pipeline_dffe[2]~q ;
wire \u19|u0|auto_generated|dffe3~q ;
wire \u20|u0|auto_generated|pipeline_dffe[3]~q ;
wire \u19|u0|auto_generated|dffe4~q ;
wire \u20|u0|auto_generated|pipeline_dffe[4]~q ;
wire \u19|u0|auto_generated|dffe5~q ;
wire \u20|u0|auto_generated|pipeline_dffe[5]~q ;
wire \u19|u0|auto_generated|dffe6~q ;
wire \u20|u0|auto_generated|pipeline_dffe[6]~q ;
wire \u19|u0|auto_generated|dffe7~q ;
wire \u24|u0|auto_generated|dffe2~q ;
wire \u21|u0|auto_generated|dffe5~q ;
wire \u18|u0|auto_generated|dffe8~q ;
wire \u15|u0|auto_generated|dffe11~q ;
wire \u12|u0|auto_generated|dffe14~q ;
wire \u9|u0|auto_generated|dffe16~q ;
wire \u16|u0|auto_generated|dffe10~q ;
wire \u14|u0|auto_generated|pipeline_dffe[12]~q ;
wire \u10|u0|auto_generated|dffe16~q ;
wire \u7|u0|auto_generated|dffe18~q ;
wire \u17|u0|auto_generated|pipeline_dffe[9]~q ;
wire \u13|u0|auto_generated|dffe13~q ;
wire \u11|u0|auto_generated|pipeline_dffe[15]~q ;
wire \u8|u0|auto_generated|pipeline_dffe[17]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[25]~q ;
wire \u24|u0|auto_generated|dffe1~q ;
wire \u21|u0|auto_generated|dffe4~q ;
wire \u18|u0|auto_generated|dffe7~q ;
wire \u15|u0|auto_generated|dffe10~q ;
wire \u12|u0|auto_generated|dffe13~q ;
wire \u16|u0|auto_generated|dffe9~q ;
wire \u14|u0|auto_generated|pipeline_dffe[11]~q ;
wire \u10|u0|auto_generated|dffe15~q ;
wire \u17|u0|auto_generated|pipeline_dffe[8]~q ;
wire \u13|u0|auto_generated|dffe12~q ;
wire \u11|u0|auto_generated|pipeline_dffe[14]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[24]~q ;
wire \u16|u0|auto_generated|dffe7~q ;
wire \u16|u0|auto_generated|dffe8~q ;
wire \u21|u0|auto_generated|dffe3~q ;
wire \u18|u0|auto_generated|dffe6~q ;
wire \u15|u0|auto_generated|dffe9~q ;
wire \u12|u0|auto_generated|dffe12~q ;
wire \u9|u0|auto_generated|dffe15~q ;
wire \u14|u0|auto_generated|pipeline_dffe[10]~q ;
wire \u10|u0|auto_generated|dffe14~q ;
wire \u8|u0|auto_generated|pipeline_dffe[16]~q ;
wire \u17|u0|auto_generated|pipeline_dffe[6]~q ;
wire \u17|u0|auto_generated|pipeline_dffe[7]~q ;
wire \u13|u0|auto_generated|dffe11~q ;
wire \u11|u0|auto_generated|pipeline_dffe[13]~q ;
wire \u7|u0|auto_generated|dffe17~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[23]~q ;
wire \u17|u0|auto_generated|pipeline_dffe[0]~q ;
wire \u21|u0|auto_generated|dffe2~q ;
wire \u18|u0|auto_generated|dffe5~q ;
wire \u15|u0|auto_generated|dffe8~q ;
wire \u12|u0|auto_generated|dffe11~q ;
wire \u9|u0|auto_generated|dffe14~q ;
wire \u6|u0|auto_generated|dffe16~q ;
wire \u14|u0|auto_generated|pipeline_dffe[9]~q ;
wire \u10|u0|auto_generated|dffe13~q ;
wire \u8|u0|auto_generated|pipeline_dffe[15]~q ;
wire \u5|u0|auto_generated|pipeline_dffe[17]~q ;
wire \u16|u0|auto_generated|dffe1~q ;
wire \u13|u0|auto_generated|dffe10~q ;
wire \u11|u0|auto_generated|pipeline_dffe[12]~q ;
wire \u7|u0|auto_generated|dffe16~q ;
wire \u4|u0|auto_generated|dffe18~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[22]~q ;
wire \u17|u0|auto_generated|pipeline_dffe[1]~q ;
wire \u16|u0|auto_generated|dffe2~q ;
wire \u17|u0|auto_generated|pipeline_dffe[2]~q ;
wire \u16|u0|auto_generated|dffe3~q ;
wire \u17|u0|auto_generated|pipeline_dffe[3]~q ;
wire \u16|u0|auto_generated|dffe4~q ;
wire \u17|u0|auto_generated|pipeline_dffe[4]~q ;
wire \u16|u0|auto_generated|dffe5~q ;
wire \u17|u0|auto_generated|pipeline_dffe[5]~q ;
wire \u16|u0|auto_generated|dffe6~q ;
wire \u21|u0|auto_generated|dffe1~q ;
wire \u18|u0|auto_generated|dffe4~q ;
wire \u15|u0|auto_generated|dffe7~q ;
wire \u12|u0|auto_generated|dffe10~q ;
wire \u9|u0|auto_generated|dffe13~q ;
wire \u14|u0|auto_generated|pipeline_dffe[8]~q ;
wire \u10|u0|auto_generated|dffe12~q ;
wire \u8|u0|auto_generated|pipeline_dffe[14]~q ;
wire \u13|u0|auto_generated|dffe9~q ;
wire \u11|u0|auto_generated|pipeline_dffe[11]~q ;
wire \u7|u0|auto_generated|dffe15~q ;
wire \u5|u0|auto_generated|pipeline_dffe[16]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[21]~q ;
wire \u18|u0|auto_generated|dffe3~q ;
wire \u15|u0|auto_generated|dffe6~q ;
wire \u12|u0|auto_generated|dffe9~q ;
wire \u9|u0|auto_generated|dffe12~q ;
wire \u6|u0|auto_generated|dffe15~q ;
wire \u14|u0|auto_generated|pipeline_dffe[7]~q ;
wire \u10|u0|auto_generated|dffe11~q ;
wire \u8|u0|auto_generated|pipeline_dffe[13]~q ;
wire \u4|u0|auto_generated|dffe17~q ;
wire \u3|u0|auto_generated|dffe16~q ;
wire \u5|xordvalue~0_combout ;
wire \u13|u0|auto_generated|dffe8~q ;
wire \u11|u0|auto_generated|pipeline_dffe[10]~q ;
wire \u7|u0|auto_generated|dffe14~q ;
wire \u5|u0|auto_generated|pipeline_dffe[15]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[20]~q ;
wire \u13|u0|auto_generated|dffe6~q ;
wire \u13|u0|auto_generated|dffe7~q ;
wire \u18|u0|auto_generated|dffe2~q ;
wire \u15|u0|auto_generated|dffe5~q ;
wire \u12|u0|auto_generated|dffe8~q ;
wire \u9|u0|auto_generated|dffe11~q ;
wire \u6|u0|auto_generated|dffe14~q ;
wire \u14|u0|auto_generated|pipeline_dffe[6]~q ;
wire \u10|u0|auto_generated|dffe10~q ;
wire \u8|u0|auto_generated|pipeline_dffe[12]~q ;
wire \u4|u0|auto_generated|dffe16~q ;
wire \ci|corx[10]~q ;
wire \u14|u0|auto_generated|pipeline_dffe[5]~q ;
wire \u11|u0|auto_generated|pipeline_dffe[9]~q ;
wire \u7|u0|auto_generated|dffe13~q ;
wire \u5|u0|auto_generated|pipeline_dffe[14]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[19]~q ;
wire \u14|u0|auto_generated|pipeline_dffe[0]~q ;
wire \u18|u0|auto_generated|dffe1~q ;
wire \u15|u0|auto_generated|dffe4~q ;
wire \u12|u0|auto_generated|dffe7~q ;
wire \u9|u0|auto_generated|dffe10~q ;
wire \u6|u0|auto_generated|dffe13~q ;
wire \u10|u0|auto_generated|dffe9~q ;
wire \u8|u0|auto_generated|pipeline_dffe[11]~q ;
wire \u4|u0|auto_generated|dffe15~q ;
wire \u13|u0|auto_generated|dffe1~q ;
wire \u11|u0|auto_generated|pipeline_dffe[8]~q ;
wire \u7|u0|auto_generated|dffe12~q ;
wire \u5|u0|auto_generated|pipeline_dffe[13]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[18]~q ;
wire \u14|u0|auto_generated|pipeline_dffe[1]~q ;
wire \u13|u0|auto_generated|dffe2~q ;
wire \u14|u0|auto_generated|pipeline_dffe[2]~q ;
wire \u13|u0|auto_generated|dffe3~q ;
wire \u14|u0|auto_generated|pipeline_dffe[3]~q ;
wire \u13|u0|auto_generated|dffe4~q ;
wire \u14|u0|auto_generated|pipeline_dffe[4]~q ;
wire \u13|u0|auto_generated|dffe5~q ;
wire \u15|u0|auto_generated|dffe3~q ;
wire \u12|u0|auto_generated|dffe6~q ;
wire \u9|u0|auto_generated|dffe9~q ;
wire \u6|u0|auto_generated|dffe12~q ;
wire \u3|u0|auto_generated|dffe15~q ;
wire \u10|u0|auto_generated|dffe8~q ;
wire \u8|u0|auto_generated|pipeline_dffe[10]~q ;
wire \u4|u0|auto_generated|dffe14~q ;
wire \u11|u0|auto_generated|pipeline_dffe[7]~q ;
wire \u7|u0|auto_generated|dffe11~q ;
wire \u5|u0|auto_generated|pipeline_dffe[12]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[17]~q ;
wire \u15|u0|auto_generated|dffe2~q ;
wire \u12|u0|auto_generated|dffe5~q ;
wire \u9|u0|auto_generated|dffe8~q ;
wire \u6|u0|auto_generated|dffe11~q ;
wire \u3|u0|auto_generated|dffe14~q ;
wire \u10|u0|auto_generated|dffe7~q ;
wire \u8|u0|auto_generated|pipeline_dffe[9]~q ;
wire \u4|u0|auto_generated|dffe13~q ;
wire \u11|u0|auto_generated|pipeline_dffe[6]~q ;
wire \u7|u0|auto_generated|dffe10~q ;
wire \u5|u0|auto_generated|pipeline_dffe[11]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[16]~q ;
wire \u10|u0|auto_generated|dffe5~q ;
wire \u10|u0|auto_generated|dffe6~q ;
wire \u15|u0|auto_generated|dffe1~q ;
wire \u12|u0|auto_generated|dffe4~q ;
wire \u9|u0|auto_generated|dffe7~q ;
wire \u6|u0|auto_generated|dffe10~q ;
wire \u3|u0|auto_generated|dffe13~q ;
wire \u8|u0|auto_generated|pipeline_dffe[8]~q ;
wire \u4|u0|auto_generated|dffe12~q ;
wire \u11|u0|auto_generated|pipeline_dffe[4]~q ;
wire \u11|u0|auto_generated|pipeline_dffe[5]~q ;
wire \u7|u0|auto_generated|dffe9~q ;
wire \u5|u0|auto_generated|pipeline_dffe[10]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[15]~q ;
wire \u11|u0|auto_generated|pipeline_dffe[0]~q ;
wire \u12|u0|auto_generated|dffe3~q ;
wire \u9|u0|auto_generated|dffe6~q ;
wire \u6|u0|auto_generated|dffe9~q ;
wire \u3|u0|auto_generated|dffe12~q ;
wire \u8|u0|auto_generated|pipeline_dffe[7]~q ;
wire \u4|u0|auto_generated|dffe11~q ;
wire \u10|u0|auto_generated|dffe1~q ;
wire \u7|u0|auto_generated|dffe8~q ;
wire \u5|u0|auto_generated|pipeline_dffe[9]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[14]~q ;
wire \u11|u0|auto_generated|pipeline_dffe[1]~q ;
wire \u10|u0|auto_generated|dffe2~q ;
wire \u11|u0|auto_generated|pipeline_dffe[2]~q ;
wire \u10|u0|auto_generated|dffe3~q ;
wire \u11|u0|auto_generated|pipeline_dffe[3]~q ;
wire \u10|u0|auto_generated|dffe4~q ;
wire \u12|u0|auto_generated|dffe2~q ;
wire \u9|u0|auto_generated|dffe5~q ;
wire \u6|u0|auto_generated|dffe8~q ;
wire \u3|u0|auto_generated|dffe11~q ;
wire \u8|u0|auto_generated|pipeline_dffe[6]~q ;
wire \u4|u0|auto_generated|dffe10~q ;
wire \u7|u0|auto_generated|dffe7~q ;
wire \u5|u0|auto_generated|pipeline_dffe[8]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[13]~q ;
wire \u12|u0|auto_generated|dffe1~q ;
wire \u9|u0|auto_generated|dffe4~q ;
wire \u6|u0|auto_generated|dffe7~q ;
wire \u3|u0|auto_generated|dffe10~q ;
wire \u8|u0|auto_generated|pipeline_dffe[5]~q ;
wire \u4|u0|auto_generated|dffe9~q ;
wire \u7|u0|auto_generated|dffe6~q ;
wire \u5|u0|auto_generated|pipeline_dffe[7]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[12]~q ;
wire \u7|u0|auto_generated|dffe4~q ;
wire \u7|u0|auto_generated|dffe5~q ;
wire \u9|u0|auto_generated|dffe3~q ;
wire \u6|u0|auto_generated|dffe6~q ;
wire \u3|u0|auto_generated|dffe9~q ;
wire \u8|u0|auto_generated|pipeline_dffe[4]~q ;
wire \u4|u0|auto_generated|dffe8~q ;
wire \u8|u0|auto_generated|pipeline_dffe[3]~q ;
wire \u5|u0|auto_generated|pipeline_dffe[6]~q ;
wire \ux000|acc|auto_generated|pipeline_dffe[11]~q ;
wire \u8|u0|auto_generated|pipeline_dffe[0]~q ;
wire \u9|u0|auto_generated|dffe2~q ;
wire \u6|u0|auto_generated|dffe5~q ;
wire \u3|u0|auto_generated|dffe8~q ;
wire \u4|u0|auto_generated|dffe7~q ;
wire \u7|u0|auto_generated|dffe1~q ;
wire \u5|u0|auto_generated|pipeline_dffe[5]~q ;
wire \u8|u0|auto_generated|pipeline_dffe[1]~q ;
wire \u7|u0|auto_generated|dffe2~q ;
wire \u8|u0|auto_generated|pipeline_dffe[2]~q ;
wire \u7|u0|auto_generated|dffe3~q ;
wire \u9|u0|auto_generated|dffe1~q ;
wire \u6|u0|auto_generated|dffe4~q ;
wire \u3|u0|auto_generated|dffe7~q ;
wire \u4|u0|auto_generated|dffe6~q ;
wire \u5|u0|auto_generated|pipeline_dffe[4]~q ;
wire \u6|u0|auto_generated|dffe3~q ;
wire \u3|u0|auto_generated|dffe6~q ;
wire \u4|u0|auto_generated|dffe5~q ;
wire \u5|u0|auto_generated|pipeline_dffe[3]~q ;
wire \u4|u0|auto_generated|dffe3~q ;
wire \u4|u0|auto_generated|dffe4~q ;
wire \u6|u0|auto_generated|dffe2~q ;
wire \u3|u0|auto_generated|dffe5~q ;
wire \u5|u0|auto_generated|pipeline_dffe[2]~q ;
wire \u5|u0|auto_generated|pipeline_dffe[1]~q ;
wire \u6|u0|auto_generated|dffe1~q ;
wire \u3|u0|auto_generated|dffe4~q ;
wire \u4|u0|auto_generated|dffe1~q ;
wire \u4|u0|auto_generated|dffe2~q ;
wire \u3|u0|auto_generated|dffe3~q ;
wire \u3|u0|auto_generated|dffe2~q ;
wire \u3|u0|auto_generated|dffe1~q ;
wire \u12|u0|auto_generated|dffe16~_wirecell_combout ;
wire \u15|u0|auto_generated|dffe16~_wirecell_combout ;
wire \u18|u0|auto_generated|dffe16~_wirecell_combout ;
wire \u21|u0|auto_generated|dffe16~_wirecell_combout ;
wire \u24|u0|auto_generated|dffe16~_wirecell_combout ;
wire \u27|u0|auto_generated|dffe16~_wirecell_combout ;
wire \u30|u0|auto_generated|dffe16~_wirecell_combout ;
wire \u33|u0|auto_generated|dffe16~_wirecell_combout ;
wire \u36|u0|auto_generated|dffe16~_wirecell_combout ;
wire \u39|u0|auto_generated|dffe16~_wirecell_combout ;
wire \u3|u0|auto_generated|dffe16~_wirecell_combout ;
wire \u42|u0|auto_generated|dffe16~_wirecell_combout ;
wire \u6|u0|auto_generated|dffe16~_wirecell_combout ;
wire \u9|u0|auto_generated|dffe16~_wirecell_combout ;


nco_test_cord_init ci(
	.corz_14(\ci|corz[14]~q ),
	.dxxpdo_18(\ux002|dxxpdo[18]~q ),
	.corz_13(\ci|corz[13]~q ),
	.dxxpdo_17(\ux002|dxxpdo[17]~q ),
	.corz_12(\ci|corz[12]~q ),
	.dxxpdo_16(\ux002|dxxpdo[16]~q ),
	.corz_11(\ci|corz[11]~q ),
	.dxxpdo_15(\ux002|dxxpdo[15]~q ),
	.corz_10(\ci|corz[10]~q ),
	.dxxpdo_14(\ux002|dxxpdo[14]~q ),
	.corz_9(\ci|corz[9]~q ),
	.dxxpdo_13(\ux002|dxxpdo[13]~q ),
	.corz_8(\ci|corz[8]~q ),
	.dxxpdo_12(\ux002|dxxpdo[12]~q ),
	.corz_7(\ci|corz[7]~q ),
	.dxxpdo_11(\ux002|dxxpdo[11]~q ),
	.corz_6(\ci|corz[6]~q ),
	.dxxpdo_10(\ux002|dxxpdo[10]~q ),
	.corz_5(\ci|corz[5]~q ),
	.dxxpdo_9(\ux002|dxxpdo[9]~q ),
	.corz_4(\ci|corz[4]~q ),
	.dxxpdo_8(\ux002|dxxpdo[8]~q ),
	.corz_3(\ci|corz[3]~q ),
	.dxxpdo_7(\ux002|dxxpdo[7]~q ),
	.corz_2(\ci|corz[2]~q ),
	.dxxpdo_6(\ux002|dxxpdo[6]~q ),
	.corz_1(\ci|corz[1]~q ),
	.dxxpdo_5(\ux002|dxxpdo[5]~q ),
	.corz_0(\ci|corz[0]~q ),
	.dxxpdo_4(\ux002|dxxpdo[4]~q ),
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.corx_10(\ci|corx[10]~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_asj_dxx ux002(
	.dxxpdo_20(\ux002|dxxpdo[20]~q ),
	.dxxpdo_19(\ux002|dxxpdo[19]~q ),
	.dxxrv_7(\ux001|dxxrv[7]~q ),
	.dxxrv_6(\ux001|dxxrv[6]~q ),
	.dxxrv_5(\ux001|dxxrv[5]~q ),
	.dxxpdo_18(\ux002|dxxpdo[18]~q ),
	.dxxrv_4(\ux001|dxxrv[4]~q ),
	.dxxpdo_17(\ux002|dxxpdo[17]~q ),
	.dxxrv_3(\ux001|dxxrv[3]~q ),
	.dxxpdo_16(\ux002|dxxpdo[16]~q ),
	.dxxrv_2(\ux001|dxxrv[2]~q ),
	.dxxpdo_15(\ux002|dxxpdo[15]~q ),
	.dxxrv_1(\ux001|dxxrv[1]~q ),
	.dxxpdo_14(\ux002|dxxpdo[14]~q ),
	.dxxrv_0(\ux001|dxxrv[0]~q ),
	.dxxpdo_13(\ux002|dxxpdo[13]~q ),
	.dxxpdo_12(\ux002|dxxpdo[12]~q ),
	.dxxpdo_11(\ux002|dxxpdo[11]~q ),
	.dxxpdo_10(\ux002|dxxpdo[10]~q ),
	.dxxpdo_9(\ux002|dxxpdo[9]~q ),
	.dxxpdo_8(\ux002|dxxpdo[8]~q ),
	.dxxpdo_7(\ux002|dxxpdo[7]~q ),
	.dxxpdo_6(\ux002|dxxpdo[6]~q ),
	.dxxpdo_5(\ux002|dxxpdo[5]~q ),
	.dxxpdo_4(\ux002|dxxpdo[4]~q ),
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.pipeline_dffe_31(\ux000|acc|auto_generated|pipeline_dffe[31]~q ),
	.pipeline_dffe_30(\ux000|acc|auto_generated|pipeline_dffe[30]~q ),
	.pipeline_dffe_29(\ux000|acc|auto_generated|pipeline_dffe[29]~q ),
	.pipeline_dffe_28(\ux000|acc|auto_generated|pipeline_dffe[28]~q ),
	.pipeline_dffe_27(\ux000|acc|auto_generated|pipeline_dffe[27]~q ),
	.pipeline_dffe_26(\ux000|acc|auto_generated|pipeline_dffe[26]~q ),
	.pipeline_dffe_25(\ux000|acc|auto_generated|pipeline_dffe[25]~q ),
	.pipeline_dffe_24(\ux000|acc|auto_generated|pipeline_dffe[24]~q ),
	.pipeline_dffe_23(\ux000|acc|auto_generated|pipeline_dffe[23]~q ),
	.pipeline_dffe_22(\ux000|acc|auto_generated|pipeline_dffe[22]~q ),
	.pipeline_dffe_21(\ux000|acc|auto_generated|pipeline_dffe[21]~q ),
	.pipeline_dffe_20(\ux000|acc|auto_generated|pipeline_dffe[20]~q ),
	.pipeline_dffe_19(\ux000|acc|auto_generated|pipeline_dffe[19]~q ),
	.pipeline_dffe_18(\ux000|acc|auto_generated|pipeline_dffe[18]~q ),
	.pipeline_dffe_17(\ux000|acc|auto_generated|pipeline_dffe[17]~q ),
	.pipeline_dffe_16(\ux000|acc|auto_generated|pipeline_dffe[16]~q ),
	.pipeline_dffe_15(\ux000|acc|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_14(\ux000|acc|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_13(\ux000|acc|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_12(\ux000|acc|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_11(\ux000|acc|auto_generated|pipeline_dffe[11]~q ),
	.clk(clk),
	.reset_n(reset_n));

nco_test_asj_dxx_g ux001(
	.dxxrv_7(\ux001|dxxrv[7]~q ),
	.dxxrv_6(\ux001|dxxrv[6]~q ),
	.dxxrv_5(\ux001|dxxrv[5]~q ),
	.dxxrv_4(\ux001|dxxrv[4]~q ),
	.dxxrv_3(\ux001|dxxrv[3]~q ),
	.dxxrv_2(\ux001|dxxrv[2]~q ),
	.dxxrv_1(\ux001|dxxrv[1]~q ),
	.dxxrv_0(\ux001|dxxrv[0]~q ),
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.clk(clk),
	.reset_n(reset_n));

nco_test_asj_altqmcpipe ux000(
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.pipeline_dffe_31(\ux000|acc|auto_generated|pipeline_dffe[31]~q ),
	.pipeline_dffe_30(\ux000|acc|auto_generated|pipeline_dffe[30]~q ),
	.pipeline_dffe_29(\ux000|acc|auto_generated|pipeline_dffe[29]~q ),
	.pipeline_dffe_28(\ux000|acc|auto_generated|pipeline_dffe[28]~q ),
	.pipeline_dffe_27(\ux000|acc|auto_generated|pipeline_dffe[27]~q ),
	.pipeline_dffe_26(\ux000|acc|auto_generated|pipeline_dffe[26]~q ),
	.pipeline_dffe_25(\ux000|acc|auto_generated|pipeline_dffe[25]~q ),
	.pipeline_dffe_24(\ux000|acc|auto_generated|pipeline_dffe[24]~q ),
	.pipeline_dffe_23(\ux000|acc|auto_generated|pipeline_dffe[23]~q ),
	.pipeline_dffe_22(\ux000|acc|auto_generated|pipeline_dffe[22]~q ),
	.pipeline_dffe_21(\ux000|acc|auto_generated|pipeline_dffe[21]~q ),
	.pipeline_dffe_20(\ux000|acc|auto_generated|pipeline_dffe[20]~q ),
	.pipeline_dffe_19(\ux000|acc|auto_generated|pipeline_dffe[19]~q ),
	.pipeline_dffe_18(\ux000|acc|auto_generated|pipeline_dffe[18]~q ),
	.pipeline_dffe_17(\ux000|acc|auto_generated|pipeline_dffe[17]~q ),
	.pipeline_dffe_16(\ux000|acc|auto_generated|pipeline_dffe[16]~q ),
	.pipeline_dffe_15(\ux000|acc|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_14(\ux000|acc|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_13(\ux000|acc|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_12(\ux000|acc|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_11(\ux000|acc|auto_generated|pipeline_dffe[11]~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken),
	.phi_inc_i_31(phi_inc_i_31),
	.phi_inc_i_30(phi_inc_i_30),
	.phi_inc_i_29(phi_inc_i_29),
	.phi_inc_i_28(phi_inc_i_28),
	.phi_inc_i_27(phi_inc_i_27),
	.phi_inc_i_26(phi_inc_i_26),
	.phi_inc_i_25(phi_inc_i_25),
	.phi_inc_i_24(phi_inc_i_24),
	.phi_inc_i_23(phi_inc_i_23),
	.phi_inc_i_22(phi_inc_i_22),
	.phi_inc_i_21(phi_inc_i_21),
	.phi_inc_i_20(phi_inc_i_20),
	.phi_inc_i_19(phi_inc_i_19),
	.phi_inc_i_18(phi_inc_i_18),
	.phi_inc_i_17(phi_inc_i_17),
	.phi_inc_i_16(phi_inc_i_16),
	.phi_inc_i_15(phi_inc_i_15),
	.phi_inc_i_14(phi_inc_i_14),
	.phi_inc_i_13(phi_inc_i_13),
	.phi_inc_i_12(phi_inc_i_12),
	.phi_inc_i_11(phi_inc_i_11),
	.phi_inc_i_10(phi_inc_i_10),
	.phi_inc_i_9(phi_inc_i_9),
	.phi_inc_i_8(phi_inc_i_8),
	.phi_inc_i_7(phi_inc_i_7),
	.phi_inc_i_6(phi_inc_i_6),
	.phi_inc_i_5(phi_inc_i_5),
	.phi_inc_i_4(phi_inc_i_4),
	.phi_inc_i_3(phi_inc_i_3),
	.phi_inc_i_2(phi_inc_i_2),
	.phi_inc_i_1(phi_inc_i_1),
	.phi_inc_i_0(phi_inc_i_0));

nco_test_cord_seg_sel css(
	.seg_rot_1(\css|seg_rot[1]~q ),
	.seg_rot_0(\css|seg_rot[0]~q ),
	.dxxpdo_20(\ux002|dxxpdo[20]~q ),
	.dxxpdo_19(\ux002|dxxpdo[19]~q ),
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.clk(clk),
	.reset_n(reset_n));

nco_test_cord_fs cfs(
	.cor1x_10(\cfs|cor1x[10]~q ),
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.corx_10(\ci|corx[10]~q ),
	.clk(clk),
	.reset_n(reset_n));

nco_test_cordic_sxor_1p_lpm_10 u4(
	.a_0(\u5|a[0]~q ),
	.xordvalue_11(\u5|xordvalue[11]~q ),
	.cor1x_10(\cfs|cor1x[10]~q ),
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.dffe18(\u4|u0|auto_generated|dffe18~q ),
	.dffe17(\u4|u0|auto_generated|dffe17~q ),
	.dffe16(\u3|u0|auto_generated|dffe16~q ),
	.xordvalue(\u5|xordvalue~0_combout ),
	.dffe161(\u4|u0|auto_generated|dffe16~q ),
	.dffe15(\u4|u0|auto_generated|dffe15~q ),
	.dffe14(\u4|u0|auto_generated|dffe14~q ),
	.dffe13(\u4|u0|auto_generated|dffe13~q ),
	.dffe12(\u4|u0|auto_generated|dffe12~q ),
	.dffe11(\u4|u0|auto_generated|dffe11~q ),
	.dffe10(\u4|u0|auto_generated|dffe10~q ),
	.dffe9(\u4|u0|auto_generated|dffe9~q ),
	.dffe8(\u4|u0|auto_generated|dffe8~q ),
	.dffe7(\u4|u0|auto_generated|dffe7~q ),
	.dffe6(\u4|u0|auto_generated|dffe6~q ),
	.dffe5(\u4|u0|auto_generated|dffe5~q ),
	.dffe3(\u4|u0|auto_generated|dffe3~q ),
	.dffe4(\u4|u0|auto_generated|dffe4~q ),
	.dffe1(\u4|u0|auto_generated|dffe1~q ),
	.dffe2(\u4|u0|auto_generated|dffe2~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_cordic_zxor_1p_lpm_6 u3(
	.corz_14(\ci|corz[14]~q ),
	.corz_13(\ci|corz[13]~q ),
	.corz_12(\ci|corz[12]~q ),
	.corz_11(\ci|corz[11]~q ),
	.corz_10(\ci|corz[10]~q ),
	.corz_9(\ci|corz[9]~q ),
	.corz_8(\ci|corz[8]~q ),
	.corz_7(\ci|corz[7]~q ),
	.corz_6(\ci|corz[6]~q ),
	.corz_5(\ci|corz[5]~q ),
	.corz_4(\ci|corz[4]~q ),
	.corz_3(\ci|corz[3]~q ),
	.corz_2(\ci|corz[2]~q ),
	.corz_1(\ci|corz[1]~q ),
	.corz_0(\ci|corz[0]~q ),
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.dffe16(\u3|u0|auto_generated|dffe16~q ),
	.corx_10(\ci|corx[10]~q ),
	.dffe15(\u3|u0|auto_generated|dffe15~q ),
	.dffe14(\u3|u0|auto_generated|dffe14~q ),
	.dffe13(\u3|u0|auto_generated|dffe13~q ),
	.dffe12(\u3|u0|auto_generated|dffe12~q ),
	.dffe11(\u3|u0|auto_generated|dffe11~q ),
	.dffe10(\u3|u0|auto_generated|dffe10~q ),
	.dffe9(\u3|u0|auto_generated|dffe9~q ),
	.dffe8(\u3|u0|auto_generated|dffe8~q ),
	.dffe7(\u3|u0|auto_generated|dffe7~q ),
	.dffe6(\u3|u0|auto_generated|dffe6~q ),
	.dffe5(\u3|u0|auto_generated|dffe5~q ),
	.dffe4(\u3|u0|auto_generated|dffe4~q ),
	.dffe3(\u3|u0|auto_generated|dffe3~q ),
	.dffe2(\u3|u0|auto_generated|dffe2~q ),
	.dffe1(\u3|u0|auto_generated|dffe1~q ),
	.dffe161(\u3|u0|auto_generated|dffe16~_wirecell_combout ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_cordic_zxor_1p_lpm_15 u6(
	.a_0(\u5|a[0]~q ),
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.dffe16(\u6|u0|auto_generated|dffe16~q ),
	.dffe15(\u6|u0|auto_generated|dffe15~q ),
	.dffe161(\u3|u0|auto_generated|dffe16~q ),
	.dffe14(\u6|u0|auto_generated|dffe14~q ),
	.dffe13(\u6|u0|auto_generated|dffe13~q ),
	.dffe12(\u6|u0|auto_generated|dffe12~q ),
	.dffe151(\u3|u0|auto_generated|dffe15~q ),
	.dffe11(\u6|u0|auto_generated|dffe11~q ),
	.dffe141(\u3|u0|auto_generated|dffe14~q ),
	.dffe10(\u6|u0|auto_generated|dffe10~q ),
	.dffe131(\u3|u0|auto_generated|dffe13~q ),
	.dffe9(\u6|u0|auto_generated|dffe9~q ),
	.dffe121(\u3|u0|auto_generated|dffe12~q ),
	.dffe8(\u6|u0|auto_generated|dffe8~q ),
	.dffe111(\u3|u0|auto_generated|dffe11~q ),
	.dffe7(\u6|u0|auto_generated|dffe7~q ),
	.dffe101(\u3|u0|auto_generated|dffe10~q ),
	.dffe6(\u6|u0|auto_generated|dffe6~q ),
	.dffe91(\u3|u0|auto_generated|dffe9~q ),
	.dffe5(\u6|u0|auto_generated|dffe5~q ),
	.dffe81(\u3|u0|auto_generated|dffe8~q ),
	.dffe4(\u6|u0|auto_generated|dffe4~q ),
	.dffe71(\u3|u0|auto_generated|dffe7~q ),
	.dffe3(\u6|u0|auto_generated|dffe3~q ),
	.dffe61(\u3|u0|auto_generated|dffe6~q ),
	.dffe2(\u6|u0|auto_generated|dffe2~q ),
	.dffe51(\u3|u0|auto_generated|dffe5~q ),
	.dffe1(\u6|u0|auto_generated|dffe1~q ),
	.dffe41(\u3|u0|auto_generated|dffe4~q ),
	.dffe31(\u3|u0|auto_generated|dffe3~q ),
	.dffe21(\u3|u0|auto_generated|dffe2~q ),
	.dffe17(\u3|u0|auto_generated|dffe1~q ),
	.dffe162(\u3|u0|auto_generated|dffe16~_wirecell_combout ),
	.dffe163(\u6|u0|auto_generated|dffe16~_wirecell_combout ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_cordic_axor_1p_lpm_13 u5(
	.a_0(\u5|a[0]~q ),
	.xordvalue_11(\u5|xordvalue[11]~q ),
	.cor1x_10(\cfs|cor1x[10]~q ),
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.pipeline_dffe_17(\u5|u0|auto_generated|pipeline_dffe[17]~q ),
	.pipeline_dffe_16(\u5|u0|auto_generated|pipeline_dffe[16]~q ),
	.dffe16(\u3|u0|auto_generated|dffe16~q ),
	.xordvalue(\u5|xordvalue~0_combout ),
	.pipeline_dffe_15(\u5|u0|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_14(\u5|u0|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_13(\u5|u0|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_12(\u5|u0|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_11(\u5|u0|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_10(\u5|u0|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_9(\u5|u0|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_8(\u5|u0|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_7(\u5|u0|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_6(\u5|u0|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_5(\u5|u0|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_4(\u5|u0|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_3(\u5|u0|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_2(\u5|u0|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_1(\u5|u0|auto_generated|pipeline_dffe[1]~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_cordic_axor_1p_lpm_16 u8(
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.pipeline_dffe_17(\u8|u0|auto_generated|pipeline_dffe[17]~q ),
	.pipeline_dffe_16(\u8|u0|auto_generated|pipeline_dffe[16]~q ),
	.dffe16(\u6|u0|auto_generated|dffe16~q ),
	.pipeline_dffe_15(\u8|u0|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_171(\u5|u0|auto_generated|pipeline_dffe[17]~q ),
	.dffe18(\u4|u0|auto_generated|dffe18~q ),
	.pipeline_dffe_14(\u8|u0|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_161(\u5|u0|auto_generated|pipeline_dffe[16]~q ),
	.pipeline_dffe_13(\u8|u0|auto_generated|pipeline_dffe[13]~q ),
	.dffe17(\u4|u0|auto_generated|dffe17~q ),
	.pipeline_dffe_151(\u5|u0|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_12(\u8|u0|auto_generated|pipeline_dffe[12]~q ),
	.dffe161(\u4|u0|auto_generated|dffe16~q ),
	.pipeline_dffe_141(\u5|u0|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_11(\u8|u0|auto_generated|pipeline_dffe[11]~q ),
	.dffe15(\u4|u0|auto_generated|dffe15~q ),
	.pipeline_dffe_131(\u5|u0|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_10(\u8|u0|auto_generated|pipeline_dffe[10]~q ),
	.dffe14(\u4|u0|auto_generated|dffe14~q ),
	.pipeline_dffe_121(\u5|u0|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_9(\u8|u0|auto_generated|pipeline_dffe[9]~q ),
	.dffe13(\u4|u0|auto_generated|dffe13~q ),
	.pipeline_dffe_111(\u5|u0|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_8(\u8|u0|auto_generated|pipeline_dffe[8]~q ),
	.dffe12(\u4|u0|auto_generated|dffe12~q ),
	.pipeline_dffe_101(\u5|u0|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_7(\u8|u0|auto_generated|pipeline_dffe[7]~q ),
	.dffe11(\u4|u0|auto_generated|dffe11~q ),
	.pipeline_dffe_91(\u5|u0|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_6(\u8|u0|auto_generated|pipeline_dffe[6]~q ),
	.dffe10(\u4|u0|auto_generated|dffe10~q ),
	.pipeline_dffe_81(\u5|u0|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_5(\u8|u0|auto_generated|pipeline_dffe[5]~q ),
	.dffe9(\u4|u0|auto_generated|dffe9~q ),
	.pipeline_dffe_71(\u5|u0|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_4(\u8|u0|auto_generated|pipeline_dffe[4]~q ),
	.dffe8(\u4|u0|auto_generated|dffe8~q ),
	.pipeline_dffe_3(\u8|u0|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_61(\u5|u0|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_0(\u8|u0|auto_generated|pipeline_dffe[0]~q ),
	.dffe7(\u4|u0|auto_generated|dffe7~q ),
	.pipeline_dffe_51(\u5|u0|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_1(\u8|u0|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_2(\u8|u0|auto_generated|pipeline_dffe[2]~q ),
	.dffe6(\u4|u0|auto_generated|dffe6~q ),
	.pipeline_dffe_41(\u5|u0|auto_generated|pipeline_dffe[4]~q ),
	.dffe5(\u4|u0|auto_generated|dffe5~q ),
	.pipeline_dffe_31(\u5|u0|auto_generated|pipeline_dffe[3]~q ),
	.dffe3(\u4|u0|auto_generated|dffe3~q ),
	.dffe4(\u4|u0|auto_generated|dffe4~q ),
	.pipeline_dffe_21(\u5|u0|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_18(\u5|u0|auto_generated|pipeline_dffe[1]~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_cordic_sxor_1p_lpm_16 u7(
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.dffe18(\u7|u0|auto_generated|dffe18~q ),
	.dffe17(\u7|u0|auto_generated|dffe17~q ),
	.dffe16(\u6|u0|auto_generated|dffe16~q ),
	.pipeline_dffe_17(\u5|u0|auto_generated|pipeline_dffe[17]~q ),
	.dffe161(\u7|u0|auto_generated|dffe16~q ),
	.dffe181(\u4|u0|auto_generated|dffe18~q ),
	.dffe15(\u7|u0|auto_generated|dffe15~q ),
	.pipeline_dffe_16(\u5|u0|auto_generated|pipeline_dffe[16]~q ),
	.dffe171(\u4|u0|auto_generated|dffe17~q ),
	.dffe14(\u7|u0|auto_generated|dffe14~q ),
	.pipeline_dffe_15(\u5|u0|auto_generated|pipeline_dffe[15]~q ),
	.dffe162(\u4|u0|auto_generated|dffe16~q ),
	.dffe13(\u7|u0|auto_generated|dffe13~q ),
	.pipeline_dffe_14(\u5|u0|auto_generated|pipeline_dffe[14]~q ),
	.dffe151(\u4|u0|auto_generated|dffe15~q ),
	.dffe12(\u7|u0|auto_generated|dffe12~q ),
	.pipeline_dffe_13(\u5|u0|auto_generated|pipeline_dffe[13]~q ),
	.dffe141(\u4|u0|auto_generated|dffe14~q ),
	.dffe11(\u7|u0|auto_generated|dffe11~q ),
	.pipeline_dffe_12(\u5|u0|auto_generated|pipeline_dffe[12]~q ),
	.dffe131(\u4|u0|auto_generated|dffe13~q ),
	.dffe10(\u7|u0|auto_generated|dffe10~q ),
	.pipeline_dffe_11(\u5|u0|auto_generated|pipeline_dffe[11]~q ),
	.dffe121(\u4|u0|auto_generated|dffe12~q ),
	.dffe9(\u7|u0|auto_generated|dffe9~q ),
	.pipeline_dffe_10(\u5|u0|auto_generated|pipeline_dffe[10]~q ),
	.dffe111(\u4|u0|auto_generated|dffe11~q ),
	.dffe8(\u7|u0|auto_generated|dffe8~q ),
	.pipeline_dffe_9(\u5|u0|auto_generated|pipeline_dffe[9]~q ),
	.dffe101(\u4|u0|auto_generated|dffe10~q ),
	.dffe7(\u7|u0|auto_generated|dffe7~q ),
	.pipeline_dffe_8(\u5|u0|auto_generated|pipeline_dffe[8]~q ),
	.dffe91(\u4|u0|auto_generated|dffe9~q ),
	.dffe6(\u7|u0|auto_generated|dffe6~q ),
	.pipeline_dffe_7(\u5|u0|auto_generated|pipeline_dffe[7]~q ),
	.dffe4(\u7|u0|auto_generated|dffe4~q ),
	.dffe5(\u7|u0|auto_generated|dffe5~q ),
	.dffe81(\u4|u0|auto_generated|dffe8~q ),
	.pipeline_dffe_6(\u5|u0|auto_generated|pipeline_dffe[6]~q ),
	.dffe71(\u4|u0|auto_generated|dffe7~q ),
	.dffe1(\u7|u0|auto_generated|dffe1~q ),
	.pipeline_dffe_5(\u5|u0|auto_generated|pipeline_dffe[5]~q ),
	.dffe2(\u7|u0|auto_generated|dffe2~q ),
	.dffe3(\u7|u0|auto_generated|dffe3~q ),
	.dffe61(\u4|u0|auto_generated|dffe6~q ),
	.pipeline_dffe_4(\u5|u0|auto_generated|pipeline_dffe[4]~q ),
	.dffe51(\u4|u0|auto_generated|dffe5~q ),
	.pipeline_dffe_3(\u5|u0|auto_generated|pipeline_dffe[3]~q ),
	.dffe31(\u4|u0|auto_generated|dffe3~q ),
	.dffe41(\u4|u0|auto_generated|dffe4~q ),
	.pipeline_dffe_2(\u5|u0|auto_generated|pipeline_dffe[2]~q ),
	.dffe19(\u4|u0|auto_generated|dffe1~q ),
	.dffe21(\u4|u0|auto_generated|dffe2~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_cordic_sxor_1p_lpm u10(
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.dffe18(\u10|u0|auto_generated|dffe18~q ),
	.dffe17(\u10|u0|auto_generated|dffe17~q ),
	.dffe16(\u9|u0|auto_generated|dffe16~q ),
	.dffe161(\u10|u0|auto_generated|dffe16~q ),
	.dffe181(\u7|u0|auto_generated|dffe18~q ),
	.pipeline_dffe_17(\u8|u0|auto_generated|pipeline_dffe[17]~q ),
	.dffe15(\u10|u0|auto_generated|dffe15~q ),
	.dffe14(\u10|u0|auto_generated|dffe14~q ),
	.pipeline_dffe_16(\u8|u0|auto_generated|pipeline_dffe[16]~q ),
	.dffe171(\u7|u0|auto_generated|dffe17~q ),
	.dffe13(\u10|u0|auto_generated|dffe13~q ),
	.pipeline_dffe_15(\u8|u0|auto_generated|pipeline_dffe[15]~q ),
	.dffe162(\u7|u0|auto_generated|dffe16~q ),
	.dffe12(\u10|u0|auto_generated|dffe12~q ),
	.pipeline_dffe_14(\u8|u0|auto_generated|pipeline_dffe[14]~q ),
	.dffe151(\u7|u0|auto_generated|dffe15~q ),
	.dffe11(\u10|u0|auto_generated|dffe11~q ),
	.pipeline_dffe_13(\u8|u0|auto_generated|pipeline_dffe[13]~q ),
	.dffe141(\u7|u0|auto_generated|dffe14~q ),
	.dffe10(\u10|u0|auto_generated|dffe10~q ),
	.pipeline_dffe_12(\u8|u0|auto_generated|pipeline_dffe[12]~q ),
	.dffe131(\u7|u0|auto_generated|dffe13~q ),
	.dffe9(\u10|u0|auto_generated|dffe9~q ),
	.pipeline_dffe_11(\u8|u0|auto_generated|pipeline_dffe[11]~q ),
	.dffe121(\u7|u0|auto_generated|dffe12~q ),
	.dffe8(\u10|u0|auto_generated|dffe8~q ),
	.pipeline_dffe_10(\u8|u0|auto_generated|pipeline_dffe[10]~q ),
	.dffe111(\u7|u0|auto_generated|dffe11~q ),
	.dffe7(\u10|u0|auto_generated|dffe7~q ),
	.pipeline_dffe_9(\u8|u0|auto_generated|pipeline_dffe[9]~q ),
	.dffe101(\u7|u0|auto_generated|dffe10~q ),
	.dffe5(\u10|u0|auto_generated|dffe5~q ),
	.dffe6(\u10|u0|auto_generated|dffe6~q ),
	.pipeline_dffe_8(\u8|u0|auto_generated|pipeline_dffe[8]~q ),
	.dffe91(\u7|u0|auto_generated|dffe9~q ),
	.pipeline_dffe_7(\u8|u0|auto_generated|pipeline_dffe[7]~q ),
	.dffe1(\u10|u0|auto_generated|dffe1~q ),
	.dffe81(\u7|u0|auto_generated|dffe8~q ),
	.dffe2(\u10|u0|auto_generated|dffe2~q ),
	.dffe3(\u10|u0|auto_generated|dffe3~q ),
	.dffe4(\u10|u0|auto_generated|dffe4~q ),
	.pipeline_dffe_6(\u8|u0|auto_generated|pipeline_dffe[6]~q ),
	.dffe71(\u7|u0|auto_generated|dffe7~q ),
	.pipeline_dffe_5(\u8|u0|auto_generated|pipeline_dffe[5]~q ),
	.dffe61(\u7|u0|auto_generated|dffe6~q ),
	.dffe41(\u7|u0|auto_generated|dffe4~q ),
	.dffe51(\u7|u0|auto_generated|dffe5~q ),
	.pipeline_dffe_4(\u8|u0|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_3(\u8|u0|auto_generated|pipeline_dffe[3]~q ),
	.dffe19(\u7|u0|auto_generated|dffe1~q ),
	.dffe21(\u7|u0|auto_generated|dffe2~q ),
	.dffe31(\u7|u0|auto_generated|dffe3~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_cordic_zxor_1p_lpm_16 u9(
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.dffe16(\u9|u0|auto_generated|dffe16~q ),
	.dffe15(\u9|u0|auto_generated|dffe15~q ),
	.dffe14(\u9|u0|auto_generated|dffe14~q ),
	.dffe161(\u6|u0|auto_generated|dffe16~q ),
	.dffe13(\u9|u0|auto_generated|dffe13~q ),
	.dffe12(\u9|u0|auto_generated|dffe12~q ),
	.dffe151(\u6|u0|auto_generated|dffe15~q ),
	.dffe11(\u9|u0|auto_generated|dffe11~q ),
	.dffe141(\u6|u0|auto_generated|dffe14~q ),
	.dffe10(\u9|u0|auto_generated|dffe10~q ),
	.dffe131(\u6|u0|auto_generated|dffe13~q ),
	.dffe9(\u9|u0|auto_generated|dffe9~q ),
	.dffe121(\u6|u0|auto_generated|dffe12~q ),
	.dffe8(\u9|u0|auto_generated|dffe8~q ),
	.dffe111(\u6|u0|auto_generated|dffe11~q ),
	.dffe7(\u9|u0|auto_generated|dffe7~q ),
	.dffe101(\u6|u0|auto_generated|dffe10~q ),
	.dffe6(\u9|u0|auto_generated|dffe6~q ),
	.dffe91(\u6|u0|auto_generated|dffe9~q ),
	.dffe5(\u9|u0|auto_generated|dffe5~q ),
	.dffe81(\u6|u0|auto_generated|dffe8~q ),
	.dffe4(\u9|u0|auto_generated|dffe4~q ),
	.dffe71(\u6|u0|auto_generated|dffe7~q ),
	.dffe3(\u9|u0|auto_generated|dffe3~q ),
	.dffe61(\u6|u0|auto_generated|dffe6~q ),
	.dffe2(\u9|u0|auto_generated|dffe2~q ),
	.dffe51(\u6|u0|auto_generated|dffe5~q ),
	.dffe1(\u9|u0|auto_generated|dffe1~q ),
	.dffe41(\u6|u0|auto_generated|dffe4~q ),
	.dffe31(\u6|u0|auto_generated|dffe3~q ),
	.dffe21(\u6|u0|auto_generated|dffe2~q ),
	.dffe17(\u6|u0|auto_generated|dffe1~q ),
	.dffe162(\u6|u0|auto_generated|dffe16~_wirecell_combout ),
	.dffe163(\u9|u0|auto_generated|dffe16~_wirecell_combout ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_cordic_zxor_1p_lpm u12(
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.dffe16(\u12|u0|auto_generated|dffe16~q ),
	.dffe15(\u12|u0|auto_generated|dffe15~q ),
	.dffe14(\u12|u0|auto_generated|dffe14~q ),
	.dffe161(\u9|u0|auto_generated|dffe16~q ),
	.dffe13(\u12|u0|auto_generated|dffe13~q ),
	.dffe12(\u12|u0|auto_generated|dffe12~q ),
	.dffe151(\u9|u0|auto_generated|dffe15~q ),
	.dffe11(\u12|u0|auto_generated|dffe11~q ),
	.dffe141(\u9|u0|auto_generated|dffe14~q ),
	.dffe10(\u12|u0|auto_generated|dffe10~q ),
	.dffe131(\u9|u0|auto_generated|dffe13~q ),
	.dffe9(\u12|u0|auto_generated|dffe9~q ),
	.dffe121(\u9|u0|auto_generated|dffe12~q ),
	.dffe8(\u12|u0|auto_generated|dffe8~q ),
	.dffe111(\u9|u0|auto_generated|dffe11~q ),
	.dffe7(\u12|u0|auto_generated|dffe7~q ),
	.dffe101(\u9|u0|auto_generated|dffe10~q ),
	.dffe6(\u12|u0|auto_generated|dffe6~q ),
	.dffe91(\u9|u0|auto_generated|dffe9~q ),
	.dffe5(\u12|u0|auto_generated|dffe5~q ),
	.dffe81(\u9|u0|auto_generated|dffe8~q ),
	.dffe4(\u12|u0|auto_generated|dffe4~q ),
	.dffe71(\u9|u0|auto_generated|dffe7~q ),
	.dffe3(\u12|u0|auto_generated|dffe3~q ),
	.dffe61(\u9|u0|auto_generated|dffe6~q ),
	.dffe2(\u12|u0|auto_generated|dffe2~q ),
	.dffe51(\u9|u0|auto_generated|dffe5~q ),
	.dffe1(\u12|u0|auto_generated|dffe1~q ),
	.dffe41(\u9|u0|auto_generated|dffe4~q ),
	.dffe31(\u9|u0|auto_generated|dffe3~q ),
	.dffe21(\u9|u0|auto_generated|dffe2~q ),
	.dffe17(\u9|u0|auto_generated|dffe1~q ),
	.dffe162(\u12|u0|auto_generated|dffe16~_wirecell_combout ),
	.dffe163(\u9|u0|auto_generated|dffe16~_wirecell_combout ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_cordic_axor_1p_lpm u11(
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.pipeline_dffe_17(\u11|u0|auto_generated|pipeline_dffe[17]~q ),
	.pipeline_dffe_16(\u11|u0|auto_generated|pipeline_dffe[16]~q ),
	.dffe16(\u9|u0|auto_generated|dffe16~q ),
	.dffe18(\u7|u0|auto_generated|dffe18~q ),
	.pipeline_dffe_15(\u11|u0|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_171(\u8|u0|auto_generated|pipeline_dffe[17]~q ),
	.pipeline_dffe_14(\u11|u0|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_161(\u8|u0|auto_generated|pipeline_dffe[16]~q ),
	.pipeline_dffe_13(\u11|u0|auto_generated|pipeline_dffe[13]~q ),
	.dffe17(\u7|u0|auto_generated|dffe17~q ),
	.pipeline_dffe_151(\u8|u0|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_12(\u11|u0|auto_generated|pipeline_dffe[12]~q ),
	.dffe161(\u7|u0|auto_generated|dffe16~q ),
	.pipeline_dffe_141(\u8|u0|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_11(\u11|u0|auto_generated|pipeline_dffe[11]~q ),
	.dffe15(\u7|u0|auto_generated|dffe15~q ),
	.pipeline_dffe_131(\u8|u0|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_10(\u11|u0|auto_generated|pipeline_dffe[10]~q ),
	.dffe14(\u7|u0|auto_generated|dffe14~q ),
	.pipeline_dffe_121(\u8|u0|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_9(\u11|u0|auto_generated|pipeline_dffe[9]~q ),
	.dffe13(\u7|u0|auto_generated|dffe13~q ),
	.pipeline_dffe_111(\u8|u0|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_8(\u11|u0|auto_generated|pipeline_dffe[8]~q ),
	.dffe12(\u7|u0|auto_generated|dffe12~q ),
	.pipeline_dffe_101(\u8|u0|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_7(\u11|u0|auto_generated|pipeline_dffe[7]~q ),
	.dffe11(\u7|u0|auto_generated|dffe11~q ),
	.pipeline_dffe_91(\u8|u0|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_6(\u11|u0|auto_generated|pipeline_dffe[6]~q ),
	.dffe10(\u7|u0|auto_generated|dffe10~q ),
	.pipeline_dffe_81(\u8|u0|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_4(\u11|u0|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\u11|u0|auto_generated|pipeline_dffe[5]~q ),
	.dffe9(\u7|u0|auto_generated|dffe9~q ),
	.pipeline_dffe_0(\u11|u0|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_71(\u8|u0|auto_generated|pipeline_dffe[7]~q ),
	.dffe8(\u7|u0|auto_generated|dffe8~q ),
	.pipeline_dffe_1(\u11|u0|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_2(\u11|u0|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\u11|u0|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_61(\u8|u0|auto_generated|pipeline_dffe[6]~q ),
	.dffe7(\u7|u0|auto_generated|dffe7~q ),
	.pipeline_dffe_51(\u8|u0|auto_generated|pipeline_dffe[5]~q ),
	.dffe6(\u7|u0|auto_generated|dffe6~q ),
	.dffe4(\u7|u0|auto_generated|dffe4~q ),
	.dffe5(\u7|u0|auto_generated|dffe5~q ),
	.pipeline_dffe_41(\u8|u0|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_31(\u8|u0|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_01(\u8|u0|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_18(\u8|u0|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_21(\u8|u0|auto_generated|pipeline_dffe[2]~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_cordic_sxor_1p_lpm_1 u13(
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.dffe18(\u13|u0|auto_generated|dffe18~q ),
	.dffe17(\u13|u0|auto_generated|dffe17~q ),
	.dffe16(\u12|u0|auto_generated|dffe16~q ),
	.pipeline_dffe_17(\u11|u0|auto_generated|pipeline_dffe[17]~q ),
	.dffe161(\u13|u0|auto_generated|dffe16~q ),
	.dffe181(\u10|u0|auto_generated|dffe18~q ),
	.dffe15(\u13|u0|auto_generated|dffe15~q ),
	.dffe171(\u10|u0|auto_generated|dffe17~q ),
	.dffe14(\u13|u0|auto_generated|dffe14~q ),
	.pipeline_dffe_16(\u11|u0|auto_generated|pipeline_dffe[16]~q ),
	.dffe162(\u10|u0|auto_generated|dffe16~q ),
	.dffe13(\u13|u0|auto_generated|dffe13~q ),
	.pipeline_dffe_15(\u11|u0|auto_generated|pipeline_dffe[15]~q ),
	.dffe151(\u10|u0|auto_generated|dffe15~q ),
	.dffe12(\u13|u0|auto_generated|dffe12~q ),
	.pipeline_dffe_14(\u11|u0|auto_generated|pipeline_dffe[14]~q ),
	.dffe141(\u10|u0|auto_generated|dffe14~q ),
	.dffe11(\u13|u0|auto_generated|dffe11~q ),
	.pipeline_dffe_13(\u11|u0|auto_generated|pipeline_dffe[13]~q ),
	.dffe131(\u10|u0|auto_generated|dffe13~q ),
	.dffe10(\u13|u0|auto_generated|dffe10~q ),
	.pipeline_dffe_12(\u11|u0|auto_generated|pipeline_dffe[12]~q ),
	.dffe121(\u10|u0|auto_generated|dffe12~q ),
	.dffe9(\u13|u0|auto_generated|dffe9~q ),
	.pipeline_dffe_11(\u11|u0|auto_generated|pipeline_dffe[11]~q ),
	.dffe111(\u10|u0|auto_generated|dffe11~q ),
	.dffe8(\u13|u0|auto_generated|dffe8~q ),
	.pipeline_dffe_10(\u11|u0|auto_generated|pipeline_dffe[10]~q ),
	.dffe6(\u13|u0|auto_generated|dffe6~q ),
	.dffe7(\u13|u0|auto_generated|dffe7~q ),
	.dffe101(\u10|u0|auto_generated|dffe10~q ),
	.pipeline_dffe_9(\u11|u0|auto_generated|pipeline_dffe[9]~q ),
	.dffe91(\u10|u0|auto_generated|dffe9~q ),
	.dffe1(\u13|u0|auto_generated|dffe1~q ),
	.pipeline_dffe_8(\u11|u0|auto_generated|pipeline_dffe[8]~q ),
	.dffe2(\u13|u0|auto_generated|dffe2~q ),
	.dffe3(\u13|u0|auto_generated|dffe3~q ),
	.dffe4(\u13|u0|auto_generated|dffe4~q ),
	.dffe5(\u13|u0|auto_generated|dffe5~q ),
	.dffe81(\u10|u0|auto_generated|dffe8~q ),
	.pipeline_dffe_7(\u11|u0|auto_generated|pipeline_dffe[7]~q ),
	.dffe71(\u10|u0|auto_generated|dffe7~q ),
	.pipeline_dffe_6(\u11|u0|auto_generated|pipeline_dffe[6]~q ),
	.dffe51(\u10|u0|auto_generated|dffe5~q ),
	.dffe61(\u10|u0|auto_generated|dffe6~q ),
	.pipeline_dffe_4(\u11|u0|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\u11|u0|auto_generated|pipeline_dffe[5]~q ),
	.dffe19(\u10|u0|auto_generated|dffe1~q ),
	.dffe21(\u10|u0|auto_generated|dffe2~q ),
	.dffe31(\u10|u0|auto_generated|dffe3~q ),
	.dffe41(\u10|u0|auto_generated|dffe4~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_cordic_zxor_1p_lpm_1 u15(
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.dffe16(\u15|u0|auto_generated|dffe16~q ),
	.dffe15(\u15|u0|auto_generated|dffe15~q ),
	.dffe14(\u15|u0|auto_generated|dffe14~q ),
	.dffe161(\u12|u0|auto_generated|dffe16~q ),
	.dffe13(\u15|u0|auto_generated|dffe13~q ),
	.dffe12(\u15|u0|auto_generated|dffe12~q ),
	.dffe151(\u12|u0|auto_generated|dffe15~q ),
	.dffe11(\u15|u0|auto_generated|dffe11~q ),
	.dffe141(\u12|u0|auto_generated|dffe14~q ),
	.dffe10(\u15|u0|auto_generated|dffe10~q ),
	.dffe131(\u12|u0|auto_generated|dffe13~q ),
	.dffe9(\u15|u0|auto_generated|dffe9~q ),
	.dffe121(\u12|u0|auto_generated|dffe12~q ),
	.dffe8(\u15|u0|auto_generated|dffe8~q ),
	.dffe111(\u12|u0|auto_generated|dffe11~q ),
	.dffe7(\u15|u0|auto_generated|dffe7~q ),
	.dffe101(\u12|u0|auto_generated|dffe10~q ),
	.dffe6(\u15|u0|auto_generated|dffe6~q ),
	.dffe91(\u12|u0|auto_generated|dffe9~q ),
	.dffe5(\u15|u0|auto_generated|dffe5~q ),
	.dffe81(\u12|u0|auto_generated|dffe8~q ),
	.dffe4(\u15|u0|auto_generated|dffe4~q ),
	.dffe71(\u12|u0|auto_generated|dffe7~q ),
	.dffe3(\u15|u0|auto_generated|dffe3~q ),
	.dffe61(\u12|u0|auto_generated|dffe6~q ),
	.dffe2(\u15|u0|auto_generated|dffe2~q ),
	.dffe51(\u12|u0|auto_generated|dffe5~q ),
	.dffe1(\u15|u0|auto_generated|dffe1~q ),
	.dffe41(\u12|u0|auto_generated|dffe4~q ),
	.dffe31(\u12|u0|auto_generated|dffe3~q ),
	.dffe21(\u12|u0|auto_generated|dffe2~q ),
	.dffe17(\u12|u0|auto_generated|dffe1~q ),
	.dffe162(\u12|u0|auto_generated|dffe16~_wirecell_combout ),
	.dffe163(\u15|u0|auto_generated|dffe16~_wirecell_combout ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_cordic_axor_1p_lpm_1 u14(
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.pipeline_dffe_17(\u14|u0|auto_generated|pipeline_dffe[17]~q ),
	.pipeline_dffe_16(\u14|u0|auto_generated|pipeline_dffe[16]~q ),
	.dffe16(\u12|u0|auto_generated|dffe16~q ),
	.pipeline_dffe_15(\u14|u0|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_171(\u11|u0|auto_generated|pipeline_dffe[17]~q ),
	.dffe18(\u10|u0|auto_generated|dffe18~q ),
	.pipeline_dffe_14(\u14|u0|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_13(\u14|u0|auto_generated|pipeline_dffe[13]~q ),
	.dffe17(\u10|u0|auto_generated|dffe17~q ),
	.pipeline_dffe_161(\u11|u0|auto_generated|pipeline_dffe[16]~q ),
	.pipeline_dffe_12(\u14|u0|auto_generated|pipeline_dffe[12]~q ),
	.dffe161(\u10|u0|auto_generated|dffe16~q ),
	.pipeline_dffe_151(\u11|u0|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_11(\u14|u0|auto_generated|pipeline_dffe[11]~q ),
	.dffe15(\u10|u0|auto_generated|dffe15~q ),
	.pipeline_dffe_141(\u11|u0|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_10(\u14|u0|auto_generated|pipeline_dffe[10]~q ),
	.dffe14(\u10|u0|auto_generated|dffe14~q ),
	.pipeline_dffe_131(\u11|u0|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_9(\u14|u0|auto_generated|pipeline_dffe[9]~q ),
	.dffe13(\u10|u0|auto_generated|dffe13~q ),
	.pipeline_dffe_121(\u11|u0|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_8(\u14|u0|auto_generated|pipeline_dffe[8]~q ),
	.dffe12(\u10|u0|auto_generated|dffe12~q ),
	.pipeline_dffe_111(\u11|u0|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_7(\u14|u0|auto_generated|pipeline_dffe[7]~q ),
	.dffe11(\u10|u0|auto_generated|dffe11~q ),
	.pipeline_dffe_101(\u11|u0|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_6(\u14|u0|auto_generated|pipeline_dffe[6]~q ),
	.dffe10(\u10|u0|auto_generated|dffe10~q ),
	.pipeline_dffe_5(\u14|u0|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_91(\u11|u0|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_0(\u14|u0|auto_generated|pipeline_dffe[0]~q ),
	.dffe9(\u10|u0|auto_generated|dffe9~q ),
	.pipeline_dffe_81(\u11|u0|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_1(\u14|u0|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_2(\u14|u0|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\u14|u0|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\u14|u0|auto_generated|pipeline_dffe[4]~q ),
	.dffe8(\u10|u0|auto_generated|dffe8~q ),
	.pipeline_dffe_71(\u11|u0|auto_generated|pipeline_dffe[7]~q ),
	.dffe7(\u10|u0|auto_generated|dffe7~q ),
	.pipeline_dffe_61(\u11|u0|auto_generated|pipeline_dffe[6]~q ),
	.dffe5(\u10|u0|auto_generated|dffe5~q ),
	.dffe6(\u10|u0|auto_generated|dffe6~q ),
	.pipeline_dffe_41(\u11|u0|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_51(\u11|u0|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_01(\u11|u0|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_18(\u11|u0|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_21(\u11|u0|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_31(\u11|u0|auto_generated|pipeline_dffe[3]~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_cordic_axor_1p_lpm_2 u17(
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.pipeline_dffe_17(\u17|u0|auto_generated|pipeline_dffe[17]~q ),
	.pipeline_dffe_16(\u17|u0|auto_generated|pipeline_dffe[16]~q ),
	.dffe16(\u15|u0|auto_generated|dffe16~q ),
	.dffe18(\u13|u0|auto_generated|dffe18~q ),
	.pipeline_dffe_15(\u17|u0|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_171(\u14|u0|auto_generated|pipeline_dffe[17]~q ),
	.pipeline_dffe_14(\u17|u0|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_161(\u14|u0|auto_generated|pipeline_dffe[16]~q ),
	.pipeline_dffe_13(\u17|u0|auto_generated|pipeline_dffe[13]~q ),
	.dffe17(\u13|u0|auto_generated|dffe17~q ),
	.pipeline_dffe_151(\u14|u0|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_12(\u17|u0|auto_generated|pipeline_dffe[12]~q ),
	.dffe161(\u13|u0|auto_generated|dffe16~q ),
	.pipeline_dffe_141(\u14|u0|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_11(\u17|u0|auto_generated|pipeline_dffe[11]~q ),
	.dffe15(\u13|u0|auto_generated|dffe15~q ),
	.pipeline_dffe_131(\u14|u0|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_10(\u17|u0|auto_generated|pipeline_dffe[10]~q ),
	.dffe14(\u13|u0|auto_generated|dffe14~q ),
	.pipeline_dffe_121(\u14|u0|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_9(\u17|u0|auto_generated|pipeline_dffe[9]~q ),
	.dffe13(\u13|u0|auto_generated|dffe13~q ),
	.pipeline_dffe_111(\u14|u0|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_8(\u17|u0|auto_generated|pipeline_dffe[8]~q ),
	.dffe12(\u13|u0|auto_generated|dffe12~q ),
	.pipeline_dffe_101(\u14|u0|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_6(\u17|u0|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\u17|u0|auto_generated|pipeline_dffe[7]~q ),
	.dffe11(\u13|u0|auto_generated|dffe11~q ),
	.pipeline_dffe_0(\u17|u0|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_91(\u14|u0|auto_generated|pipeline_dffe[9]~q ),
	.dffe10(\u13|u0|auto_generated|dffe10~q ),
	.pipeline_dffe_1(\u17|u0|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_2(\u17|u0|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\u17|u0|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\u17|u0|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\u17|u0|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_81(\u14|u0|auto_generated|pipeline_dffe[8]~q ),
	.dffe9(\u13|u0|auto_generated|dffe9~q ),
	.pipeline_dffe_71(\u14|u0|auto_generated|pipeline_dffe[7]~q ),
	.dffe8(\u13|u0|auto_generated|dffe8~q ),
	.dffe6(\u13|u0|auto_generated|dffe6~q ),
	.dffe7(\u13|u0|auto_generated|dffe7~q ),
	.pipeline_dffe_61(\u14|u0|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_51(\u14|u0|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_01(\u14|u0|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_18(\u14|u0|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_21(\u14|u0|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_31(\u14|u0|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_41(\u14|u0|auto_generated|pipeline_dffe[4]~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_cordic_sxor_1p_lpm_2 u16(
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.dffe18(\u16|u0|auto_generated|dffe18~q ),
	.dffe17(\u16|u0|auto_generated|dffe17~q ),
	.dffe16(\u15|u0|auto_generated|dffe16~q ),
	.dffe161(\u16|u0|auto_generated|dffe16~q ),
	.dffe181(\u13|u0|auto_generated|dffe18~q ),
	.pipeline_dffe_17(\u14|u0|auto_generated|pipeline_dffe[17]~q ),
	.dffe15(\u16|u0|auto_generated|dffe15~q ),
	.dffe14(\u16|u0|auto_generated|dffe14~q ),
	.pipeline_dffe_16(\u14|u0|auto_generated|pipeline_dffe[16]~q ),
	.dffe171(\u13|u0|auto_generated|dffe17~q ),
	.dffe13(\u16|u0|auto_generated|dffe13~q ),
	.pipeline_dffe_15(\u14|u0|auto_generated|pipeline_dffe[15]~q ),
	.dffe162(\u13|u0|auto_generated|dffe16~q ),
	.dffe12(\u16|u0|auto_generated|dffe12~q ),
	.pipeline_dffe_14(\u14|u0|auto_generated|pipeline_dffe[14]~q ),
	.dffe151(\u13|u0|auto_generated|dffe15~q ),
	.dffe11(\u16|u0|auto_generated|dffe11~q ),
	.pipeline_dffe_13(\u14|u0|auto_generated|pipeline_dffe[13]~q ),
	.dffe141(\u13|u0|auto_generated|dffe14~q ),
	.dffe10(\u16|u0|auto_generated|dffe10~q ),
	.pipeline_dffe_12(\u14|u0|auto_generated|pipeline_dffe[12]~q ),
	.dffe131(\u13|u0|auto_generated|dffe13~q ),
	.dffe9(\u16|u0|auto_generated|dffe9~q ),
	.pipeline_dffe_11(\u14|u0|auto_generated|pipeline_dffe[11]~q ),
	.dffe121(\u13|u0|auto_generated|dffe12~q ),
	.dffe7(\u16|u0|auto_generated|dffe7~q ),
	.dffe8(\u16|u0|auto_generated|dffe8~q ),
	.pipeline_dffe_10(\u14|u0|auto_generated|pipeline_dffe[10]~q ),
	.dffe111(\u13|u0|auto_generated|dffe11~q ),
	.pipeline_dffe_9(\u14|u0|auto_generated|pipeline_dffe[9]~q ),
	.dffe1(\u16|u0|auto_generated|dffe1~q ),
	.dffe101(\u13|u0|auto_generated|dffe10~q ),
	.dffe2(\u16|u0|auto_generated|dffe2~q ),
	.dffe3(\u16|u0|auto_generated|dffe3~q ),
	.dffe4(\u16|u0|auto_generated|dffe4~q ),
	.dffe5(\u16|u0|auto_generated|dffe5~q ),
	.dffe6(\u16|u0|auto_generated|dffe6~q ),
	.pipeline_dffe_8(\u14|u0|auto_generated|pipeline_dffe[8]~q ),
	.dffe91(\u13|u0|auto_generated|dffe9~q ),
	.pipeline_dffe_7(\u14|u0|auto_generated|pipeline_dffe[7]~q ),
	.dffe81(\u13|u0|auto_generated|dffe8~q ),
	.dffe61(\u13|u0|auto_generated|dffe6~q ),
	.dffe71(\u13|u0|auto_generated|dffe7~q ),
	.pipeline_dffe_6(\u14|u0|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_5(\u14|u0|auto_generated|pipeline_dffe[5]~q ),
	.dffe19(\u13|u0|auto_generated|dffe1~q ),
	.dffe21(\u13|u0|auto_generated|dffe2~q ),
	.dffe31(\u13|u0|auto_generated|dffe3~q ),
	.dffe41(\u13|u0|auto_generated|dffe4~q ),
	.dffe51(\u13|u0|auto_generated|dffe5~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_cordic_sxor_1p_lpm_3 u19(
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.dffe18(\u19|u0|auto_generated|dffe18~q ),
	.dffe17(\u19|u0|auto_generated|dffe17~q ),
	.dffe16(\u18|u0|auto_generated|dffe16~q ),
	.pipeline_dffe_17(\u17|u0|auto_generated|pipeline_dffe[17]~q ),
	.dffe161(\u19|u0|auto_generated|dffe16~q ),
	.dffe181(\u16|u0|auto_generated|dffe18~q ),
	.dffe15(\u19|u0|auto_generated|dffe15~q ),
	.dffe171(\u16|u0|auto_generated|dffe17~q ),
	.dffe14(\u19|u0|auto_generated|dffe14~q ),
	.pipeline_dffe_16(\u17|u0|auto_generated|pipeline_dffe[16]~q ),
	.dffe162(\u16|u0|auto_generated|dffe16~q ),
	.dffe13(\u19|u0|auto_generated|dffe13~q ),
	.pipeline_dffe_15(\u17|u0|auto_generated|pipeline_dffe[15]~q ),
	.dffe151(\u16|u0|auto_generated|dffe15~q ),
	.dffe12(\u19|u0|auto_generated|dffe12~q ),
	.pipeline_dffe_14(\u17|u0|auto_generated|pipeline_dffe[14]~q ),
	.dffe141(\u16|u0|auto_generated|dffe14~q ),
	.dffe11(\u19|u0|auto_generated|dffe11~q ),
	.pipeline_dffe_13(\u17|u0|auto_generated|pipeline_dffe[13]~q ),
	.dffe131(\u16|u0|auto_generated|dffe13~q ),
	.dffe10(\u19|u0|auto_generated|dffe10~q ),
	.pipeline_dffe_12(\u17|u0|auto_generated|pipeline_dffe[12]~q ),
	.dffe8(\u19|u0|auto_generated|dffe8~q ),
	.dffe9(\u19|u0|auto_generated|dffe9~q ),
	.dffe121(\u16|u0|auto_generated|dffe12~q ),
	.pipeline_dffe_11(\u17|u0|auto_generated|pipeline_dffe[11]~q ),
	.dffe111(\u16|u0|auto_generated|dffe11~q ),
	.dffe1(\u19|u0|auto_generated|dffe1~q ),
	.pipeline_dffe_10(\u17|u0|auto_generated|pipeline_dffe[10]~q ),
	.dffe2(\u19|u0|auto_generated|dffe2~q ),
	.dffe3(\u19|u0|auto_generated|dffe3~q ),
	.dffe4(\u19|u0|auto_generated|dffe4~q ),
	.dffe5(\u19|u0|auto_generated|dffe5~q ),
	.dffe6(\u19|u0|auto_generated|dffe6~q ),
	.dffe7(\u19|u0|auto_generated|dffe7~q ),
	.dffe101(\u16|u0|auto_generated|dffe10~q ),
	.pipeline_dffe_9(\u17|u0|auto_generated|pipeline_dffe[9]~q ),
	.dffe91(\u16|u0|auto_generated|dffe9~q ),
	.pipeline_dffe_8(\u17|u0|auto_generated|pipeline_dffe[8]~q ),
	.dffe71(\u16|u0|auto_generated|dffe7~q ),
	.dffe81(\u16|u0|auto_generated|dffe8~q ),
	.pipeline_dffe_6(\u17|u0|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\u17|u0|auto_generated|pipeline_dffe[7]~q ),
	.dffe19(\u16|u0|auto_generated|dffe1~q ),
	.dffe21(\u16|u0|auto_generated|dffe2~q ),
	.dffe31(\u16|u0|auto_generated|dffe3~q ),
	.dffe41(\u16|u0|auto_generated|dffe4~q ),
	.dffe51(\u16|u0|auto_generated|dffe5~q ),
	.dffe61(\u16|u0|auto_generated|dffe6~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_cordic_zxor_1p_lpm_2 u18(
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.dffe16(\u18|u0|auto_generated|dffe16~q ),
	.dffe15(\u18|u0|auto_generated|dffe15~q ),
	.dffe14(\u18|u0|auto_generated|dffe14~q ),
	.dffe161(\u15|u0|auto_generated|dffe16~q ),
	.dffe13(\u18|u0|auto_generated|dffe13~q ),
	.dffe12(\u18|u0|auto_generated|dffe12~q ),
	.dffe151(\u15|u0|auto_generated|dffe15~q ),
	.dffe11(\u18|u0|auto_generated|dffe11~q ),
	.dffe141(\u15|u0|auto_generated|dffe14~q ),
	.dffe10(\u18|u0|auto_generated|dffe10~q ),
	.dffe131(\u15|u0|auto_generated|dffe13~q ),
	.dffe9(\u18|u0|auto_generated|dffe9~q ),
	.dffe121(\u15|u0|auto_generated|dffe12~q ),
	.dffe8(\u18|u0|auto_generated|dffe8~q ),
	.dffe111(\u15|u0|auto_generated|dffe11~q ),
	.dffe7(\u18|u0|auto_generated|dffe7~q ),
	.dffe101(\u15|u0|auto_generated|dffe10~q ),
	.dffe6(\u18|u0|auto_generated|dffe6~q ),
	.dffe91(\u15|u0|auto_generated|dffe9~q ),
	.dffe5(\u18|u0|auto_generated|dffe5~q ),
	.dffe81(\u15|u0|auto_generated|dffe8~q ),
	.dffe4(\u18|u0|auto_generated|dffe4~q ),
	.dffe71(\u15|u0|auto_generated|dffe7~q ),
	.dffe3(\u18|u0|auto_generated|dffe3~q ),
	.dffe61(\u15|u0|auto_generated|dffe6~q ),
	.dffe2(\u18|u0|auto_generated|dffe2~q ),
	.dffe51(\u15|u0|auto_generated|dffe5~q ),
	.dffe1(\u18|u0|auto_generated|dffe1~q ),
	.dffe41(\u15|u0|auto_generated|dffe4~q ),
	.dffe31(\u15|u0|auto_generated|dffe3~q ),
	.dffe21(\u15|u0|auto_generated|dffe2~q ),
	.dffe17(\u15|u0|auto_generated|dffe1~q ),
	.dffe162(\u15|u0|auto_generated|dffe16~_wirecell_combout ),
	.dffe163(\u18|u0|auto_generated|dffe16~_wirecell_combout ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_cordic_zxor_1p_lpm_3 u21(
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.dffe16(\u21|u0|auto_generated|dffe16~q ),
	.dffe15(\u21|u0|auto_generated|dffe15~q ),
	.dffe14(\u21|u0|auto_generated|dffe14~q ),
	.dffe161(\u18|u0|auto_generated|dffe16~q ),
	.dffe13(\u21|u0|auto_generated|dffe13~q ),
	.dffe12(\u21|u0|auto_generated|dffe12~q ),
	.dffe151(\u18|u0|auto_generated|dffe15~q ),
	.dffe11(\u21|u0|auto_generated|dffe11~q ),
	.dffe141(\u18|u0|auto_generated|dffe14~q ),
	.dffe10(\u21|u0|auto_generated|dffe10~q ),
	.dffe131(\u18|u0|auto_generated|dffe13~q ),
	.dffe9(\u21|u0|auto_generated|dffe9~q ),
	.dffe121(\u18|u0|auto_generated|dffe12~q ),
	.dffe8(\u21|u0|auto_generated|dffe8~q ),
	.dffe111(\u18|u0|auto_generated|dffe11~q ),
	.dffe7(\u21|u0|auto_generated|dffe7~q ),
	.dffe101(\u18|u0|auto_generated|dffe10~q ),
	.dffe6(\u21|u0|auto_generated|dffe6~q ),
	.dffe91(\u18|u0|auto_generated|dffe9~q ),
	.dffe5(\u21|u0|auto_generated|dffe5~q ),
	.dffe81(\u18|u0|auto_generated|dffe8~q ),
	.dffe4(\u21|u0|auto_generated|dffe4~q ),
	.dffe71(\u18|u0|auto_generated|dffe7~q ),
	.dffe3(\u21|u0|auto_generated|dffe3~q ),
	.dffe61(\u18|u0|auto_generated|dffe6~q ),
	.dffe2(\u21|u0|auto_generated|dffe2~q ),
	.dffe51(\u18|u0|auto_generated|dffe5~q ),
	.dffe1(\u21|u0|auto_generated|dffe1~q ),
	.dffe41(\u18|u0|auto_generated|dffe4~q ),
	.dffe31(\u18|u0|auto_generated|dffe3~q ),
	.dffe21(\u18|u0|auto_generated|dffe2~q ),
	.dffe17(\u18|u0|auto_generated|dffe1~q ),
	.dffe162(\u18|u0|auto_generated|dffe16~_wirecell_combout ),
	.dffe163(\u21|u0|auto_generated|dffe16~_wirecell_combout ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_cordic_axor_1p_lpm_3 u20(
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.pipeline_dffe_17(\u20|u0|auto_generated|pipeline_dffe[17]~q ),
	.pipeline_dffe_16(\u20|u0|auto_generated|pipeline_dffe[16]~q ),
	.dffe16(\u18|u0|auto_generated|dffe16~q ),
	.pipeline_dffe_15(\u20|u0|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_171(\u17|u0|auto_generated|pipeline_dffe[17]~q ),
	.dffe18(\u16|u0|auto_generated|dffe18~q ),
	.pipeline_dffe_14(\u20|u0|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_13(\u20|u0|auto_generated|pipeline_dffe[13]~q ),
	.dffe17(\u16|u0|auto_generated|dffe17~q ),
	.pipeline_dffe_161(\u17|u0|auto_generated|pipeline_dffe[16]~q ),
	.pipeline_dffe_12(\u20|u0|auto_generated|pipeline_dffe[12]~q ),
	.dffe161(\u16|u0|auto_generated|dffe16~q ),
	.pipeline_dffe_151(\u17|u0|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_11(\u20|u0|auto_generated|pipeline_dffe[11]~q ),
	.dffe15(\u16|u0|auto_generated|dffe15~q ),
	.pipeline_dffe_141(\u17|u0|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_10(\u20|u0|auto_generated|pipeline_dffe[10]~q ),
	.dffe14(\u16|u0|auto_generated|dffe14~q ),
	.pipeline_dffe_131(\u17|u0|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_9(\u20|u0|auto_generated|pipeline_dffe[9]~q ),
	.dffe13(\u16|u0|auto_generated|dffe13~q ),
	.pipeline_dffe_121(\u17|u0|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_8(\u20|u0|auto_generated|pipeline_dffe[8]~q ),
	.dffe12(\u16|u0|auto_generated|dffe12~q ),
	.pipeline_dffe_7(\u20|u0|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_111(\u17|u0|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_0(\u20|u0|auto_generated|pipeline_dffe[0]~q ),
	.dffe11(\u16|u0|auto_generated|dffe11~q ),
	.pipeline_dffe_101(\u17|u0|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_1(\u20|u0|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_2(\u20|u0|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\u20|u0|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\u20|u0|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\u20|u0|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\u20|u0|auto_generated|pipeline_dffe[6]~q ),
	.dffe10(\u16|u0|auto_generated|dffe10~q ),
	.pipeline_dffe_91(\u17|u0|auto_generated|pipeline_dffe[9]~q ),
	.dffe9(\u16|u0|auto_generated|dffe9~q ),
	.pipeline_dffe_81(\u17|u0|auto_generated|pipeline_dffe[8]~q ),
	.dffe7(\u16|u0|auto_generated|dffe7~q ),
	.dffe8(\u16|u0|auto_generated|dffe8~q ),
	.pipeline_dffe_61(\u17|u0|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_71(\u17|u0|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_01(\u17|u0|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_18(\u17|u0|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_21(\u17|u0|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_31(\u17|u0|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_41(\u17|u0|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_51(\u17|u0|auto_generated|pipeline_dffe[5]~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_cordic_axor_1p_lpm_4 u23(
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.pipeline_dffe_17(\u23|u0|auto_generated|pipeline_dffe[17]~q ),
	.pipeline_dffe_16(\u23|u0|auto_generated|pipeline_dffe[16]~q ),
	.dffe16(\u21|u0|auto_generated|dffe16~q ),
	.dffe18(\u19|u0|auto_generated|dffe18~q ),
	.pipeline_dffe_15(\u23|u0|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_171(\u20|u0|auto_generated|pipeline_dffe[17]~q ),
	.pipeline_dffe_14(\u23|u0|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_161(\u20|u0|auto_generated|pipeline_dffe[16]~q ),
	.pipeline_dffe_13(\u23|u0|auto_generated|pipeline_dffe[13]~q ),
	.dffe17(\u19|u0|auto_generated|dffe17~q ),
	.pipeline_dffe_151(\u20|u0|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_12(\u23|u0|auto_generated|pipeline_dffe[12]~q ),
	.dffe161(\u19|u0|auto_generated|dffe16~q ),
	.pipeline_dffe_141(\u20|u0|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_11(\u23|u0|auto_generated|pipeline_dffe[11]~q ),
	.dffe15(\u19|u0|auto_generated|dffe15~q ),
	.pipeline_dffe_131(\u20|u0|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_10(\u23|u0|auto_generated|pipeline_dffe[10]~q ),
	.dffe14(\u19|u0|auto_generated|dffe14~q ),
	.pipeline_dffe_121(\u20|u0|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_8(\u23|u0|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\u23|u0|auto_generated|pipeline_dffe[9]~q ),
	.dffe13(\u19|u0|auto_generated|dffe13~q ),
	.pipeline_dffe_0(\u23|u0|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_111(\u20|u0|auto_generated|pipeline_dffe[11]~q ),
	.dffe12(\u19|u0|auto_generated|dffe12~q ),
	.pipeline_dffe_1(\u23|u0|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_2(\u23|u0|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\u23|u0|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\u23|u0|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\u23|u0|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\u23|u0|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\u23|u0|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_101(\u20|u0|auto_generated|pipeline_dffe[10]~q ),
	.dffe11(\u19|u0|auto_generated|dffe11~q ),
	.pipeline_dffe_91(\u20|u0|auto_generated|pipeline_dffe[9]~q ),
	.dffe10(\u19|u0|auto_generated|dffe10~q ),
	.dffe8(\u19|u0|auto_generated|dffe8~q ),
	.dffe9(\u19|u0|auto_generated|dffe9~q ),
	.pipeline_dffe_81(\u20|u0|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_71(\u20|u0|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_01(\u20|u0|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_18(\u20|u0|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_21(\u20|u0|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_31(\u20|u0|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_41(\u20|u0|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_51(\u20|u0|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_61(\u20|u0|auto_generated|pipeline_dffe[6]~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_cordic_sxor_1p_lpm_4 u22(
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.dffe18(\u22|u0|auto_generated|dffe18~q ),
	.dffe17(\u22|u0|auto_generated|dffe17~q ),
	.dffe16(\u21|u0|auto_generated|dffe16~q ),
	.dffe161(\u22|u0|auto_generated|dffe16~q ),
	.dffe181(\u19|u0|auto_generated|dffe18~q ),
	.pipeline_dffe_17(\u20|u0|auto_generated|pipeline_dffe[17]~q ),
	.dffe15(\u22|u0|auto_generated|dffe15~q ),
	.dffe14(\u22|u0|auto_generated|dffe14~q ),
	.pipeline_dffe_16(\u20|u0|auto_generated|pipeline_dffe[16]~q ),
	.dffe171(\u19|u0|auto_generated|dffe17~q ),
	.dffe13(\u22|u0|auto_generated|dffe13~q ),
	.pipeline_dffe_15(\u20|u0|auto_generated|pipeline_dffe[15]~q ),
	.dffe162(\u19|u0|auto_generated|dffe16~q ),
	.dffe12(\u22|u0|auto_generated|dffe12~q ),
	.pipeline_dffe_14(\u20|u0|auto_generated|pipeline_dffe[14]~q ),
	.dffe151(\u19|u0|auto_generated|dffe15~q ),
	.dffe11(\u22|u0|auto_generated|dffe11~q ),
	.pipeline_dffe_13(\u20|u0|auto_generated|pipeline_dffe[13]~q ),
	.dffe141(\u19|u0|auto_generated|dffe14~q ),
	.dffe9(\u22|u0|auto_generated|dffe9~q ),
	.dffe10(\u22|u0|auto_generated|dffe10~q ),
	.pipeline_dffe_12(\u20|u0|auto_generated|pipeline_dffe[12]~q ),
	.dffe131(\u19|u0|auto_generated|dffe13~q ),
	.pipeline_dffe_11(\u20|u0|auto_generated|pipeline_dffe[11]~q ),
	.dffe1(\u22|u0|auto_generated|dffe1~q ),
	.dffe121(\u19|u0|auto_generated|dffe12~q ),
	.dffe2(\u22|u0|auto_generated|dffe2~q ),
	.dffe3(\u22|u0|auto_generated|dffe3~q ),
	.dffe4(\u22|u0|auto_generated|dffe4~q ),
	.dffe5(\u22|u0|auto_generated|dffe5~q ),
	.dffe6(\u22|u0|auto_generated|dffe6~q ),
	.dffe7(\u22|u0|auto_generated|dffe7~q ),
	.dffe8(\u22|u0|auto_generated|dffe8~q ),
	.pipeline_dffe_10(\u20|u0|auto_generated|pipeline_dffe[10]~q ),
	.dffe111(\u19|u0|auto_generated|dffe11~q ),
	.pipeline_dffe_9(\u20|u0|auto_generated|pipeline_dffe[9]~q ),
	.dffe101(\u19|u0|auto_generated|dffe10~q ),
	.dffe81(\u19|u0|auto_generated|dffe8~q ),
	.dffe91(\u19|u0|auto_generated|dffe9~q ),
	.pipeline_dffe_8(\u20|u0|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_7(\u20|u0|auto_generated|pipeline_dffe[7]~q ),
	.dffe19(\u19|u0|auto_generated|dffe1~q ),
	.dffe21(\u19|u0|auto_generated|dffe2~q ),
	.dffe31(\u19|u0|auto_generated|dffe3~q ),
	.dffe41(\u19|u0|auto_generated|dffe4~q ),
	.dffe51(\u19|u0|auto_generated|dffe5~q ),
	.dffe61(\u19|u0|auto_generated|dffe6~q ),
	.dffe71(\u19|u0|auto_generated|dffe7~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_cordic_sxor_1p_lpm_5 u25(
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.dffe18(\u25|u0|auto_generated|dffe18~q ),
	.dffe17(\u25|u0|auto_generated|dffe17~q ),
	.dffe16(\u24|u0|auto_generated|dffe16~q ),
	.pipeline_dffe_17(\u23|u0|auto_generated|pipeline_dffe[17]~q ),
	.dffe161(\u25|u0|auto_generated|dffe16~q ),
	.dffe181(\u22|u0|auto_generated|dffe18~q ),
	.dffe15(\u25|u0|auto_generated|dffe15~q ),
	.dffe171(\u22|u0|auto_generated|dffe17~q ),
	.dffe14(\u25|u0|auto_generated|dffe14~q ),
	.pipeline_dffe_16(\u23|u0|auto_generated|pipeline_dffe[16]~q ),
	.dffe162(\u22|u0|auto_generated|dffe16~q ),
	.dffe13(\u25|u0|auto_generated|dffe13~q ),
	.pipeline_dffe_15(\u23|u0|auto_generated|pipeline_dffe[15]~q ),
	.dffe151(\u22|u0|auto_generated|dffe15~q ),
	.dffe12(\u25|u0|auto_generated|dffe12~q ),
	.pipeline_dffe_14(\u23|u0|auto_generated|pipeline_dffe[14]~q ),
	.dffe10(\u25|u0|auto_generated|dffe10~q ),
	.dffe11(\u25|u0|auto_generated|dffe11~q ),
	.dffe141(\u22|u0|auto_generated|dffe14~q ),
	.pipeline_dffe_13(\u23|u0|auto_generated|pipeline_dffe[13]~q ),
	.dffe131(\u22|u0|auto_generated|dffe13~q ),
	.dffe1(\u25|u0|auto_generated|dffe1~q ),
	.pipeline_dffe_12(\u23|u0|auto_generated|pipeline_dffe[12]~q ),
	.dffe2(\u25|u0|auto_generated|dffe2~q ),
	.dffe3(\u25|u0|auto_generated|dffe3~q ),
	.dffe4(\u25|u0|auto_generated|dffe4~q ),
	.dffe5(\u25|u0|auto_generated|dffe5~q ),
	.dffe6(\u25|u0|auto_generated|dffe6~q ),
	.dffe7(\u25|u0|auto_generated|dffe7~q ),
	.dffe8(\u25|u0|auto_generated|dffe8~q ),
	.dffe9(\u25|u0|auto_generated|dffe9~q ),
	.dffe121(\u22|u0|auto_generated|dffe12~q ),
	.pipeline_dffe_11(\u23|u0|auto_generated|pipeline_dffe[11]~q ),
	.dffe111(\u22|u0|auto_generated|dffe11~q ),
	.pipeline_dffe_10(\u23|u0|auto_generated|pipeline_dffe[10]~q ),
	.dffe91(\u22|u0|auto_generated|dffe9~q ),
	.dffe101(\u22|u0|auto_generated|dffe10~q ),
	.pipeline_dffe_8(\u23|u0|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\u23|u0|auto_generated|pipeline_dffe[9]~q ),
	.dffe19(\u22|u0|auto_generated|dffe1~q ),
	.dffe21(\u22|u0|auto_generated|dffe2~q ),
	.dffe31(\u22|u0|auto_generated|dffe3~q ),
	.dffe41(\u22|u0|auto_generated|dffe4~q ),
	.dffe51(\u22|u0|auto_generated|dffe5~q ),
	.dffe61(\u22|u0|auto_generated|dffe6~q ),
	.dffe71(\u22|u0|auto_generated|dffe7~q ),
	.dffe81(\u22|u0|auto_generated|dffe8~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_cordic_zxor_1p_lpm_4 u24(
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.dffe16(\u24|u0|auto_generated|dffe16~q ),
	.dffe15(\u24|u0|auto_generated|dffe15~q ),
	.dffe14(\u24|u0|auto_generated|dffe14~q ),
	.dffe161(\u21|u0|auto_generated|dffe16~q ),
	.dffe13(\u24|u0|auto_generated|dffe13~q ),
	.dffe12(\u24|u0|auto_generated|dffe12~q ),
	.dffe151(\u21|u0|auto_generated|dffe15~q ),
	.dffe11(\u24|u0|auto_generated|dffe11~q ),
	.dffe141(\u21|u0|auto_generated|dffe14~q ),
	.dffe10(\u24|u0|auto_generated|dffe10~q ),
	.dffe131(\u21|u0|auto_generated|dffe13~q ),
	.dffe9(\u24|u0|auto_generated|dffe9~q ),
	.dffe121(\u21|u0|auto_generated|dffe12~q ),
	.dffe8(\u24|u0|auto_generated|dffe8~q ),
	.dffe111(\u21|u0|auto_generated|dffe11~q ),
	.dffe7(\u24|u0|auto_generated|dffe7~q ),
	.dffe101(\u21|u0|auto_generated|dffe10~q ),
	.dffe6(\u24|u0|auto_generated|dffe6~q ),
	.dffe91(\u21|u0|auto_generated|dffe9~q ),
	.dffe5(\u24|u0|auto_generated|dffe5~q ),
	.dffe81(\u21|u0|auto_generated|dffe8~q ),
	.dffe4(\u24|u0|auto_generated|dffe4~q ),
	.dffe71(\u21|u0|auto_generated|dffe7~q ),
	.dffe3(\u24|u0|auto_generated|dffe3~q ),
	.dffe61(\u21|u0|auto_generated|dffe6~q ),
	.dffe2(\u24|u0|auto_generated|dffe2~q ),
	.dffe51(\u21|u0|auto_generated|dffe5~q ),
	.dffe1(\u24|u0|auto_generated|dffe1~q ),
	.dffe41(\u21|u0|auto_generated|dffe4~q ),
	.dffe31(\u21|u0|auto_generated|dffe3~q ),
	.dffe21(\u21|u0|auto_generated|dffe2~q ),
	.dffe17(\u21|u0|auto_generated|dffe1~q ),
	.dffe162(\u21|u0|auto_generated|dffe16~_wirecell_combout ),
	.dffe163(\u24|u0|auto_generated|dffe16~_wirecell_combout ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_cordic_zxor_1p_lpm_5 u27(
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.dffe16(\u27|u0|auto_generated|dffe16~q ),
	.dffe15(\u27|u0|auto_generated|dffe15~q ),
	.dffe14(\u27|u0|auto_generated|dffe14~q ),
	.dffe161(\u24|u0|auto_generated|dffe16~q ),
	.dffe13(\u27|u0|auto_generated|dffe13~q ),
	.dffe12(\u27|u0|auto_generated|dffe12~q ),
	.dffe151(\u24|u0|auto_generated|dffe15~q ),
	.dffe11(\u27|u0|auto_generated|dffe11~q ),
	.dffe141(\u24|u0|auto_generated|dffe14~q ),
	.dffe10(\u27|u0|auto_generated|dffe10~q ),
	.dffe131(\u24|u0|auto_generated|dffe13~q ),
	.dffe9(\u27|u0|auto_generated|dffe9~q ),
	.dffe121(\u24|u0|auto_generated|dffe12~q ),
	.dffe8(\u27|u0|auto_generated|dffe8~q ),
	.dffe111(\u24|u0|auto_generated|dffe11~q ),
	.dffe7(\u27|u0|auto_generated|dffe7~q ),
	.dffe101(\u24|u0|auto_generated|dffe10~q ),
	.dffe6(\u27|u0|auto_generated|dffe6~q ),
	.dffe91(\u24|u0|auto_generated|dffe9~q ),
	.dffe5(\u27|u0|auto_generated|dffe5~q ),
	.dffe81(\u24|u0|auto_generated|dffe8~q ),
	.dffe4(\u27|u0|auto_generated|dffe4~q ),
	.dffe71(\u24|u0|auto_generated|dffe7~q ),
	.dffe3(\u27|u0|auto_generated|dffe3~q ),
	.dffe61(\u24|u0|auto_generated|dffe6~q ),
	.dffe2(\u27|u0|auto_generated|dffe2~q ),
	.dffe51(\u24|u0|auto_generated|dffe5~q ),
	.dffe1(\u27|u0|auto_generated|dffe1~q ),
	.dffe41(\u24|u0|auto_generated|dffe4~q ),
	.dffe31(\u24|u0|auto_generated|dffe3~q ),
	.dffe21(\u24|u0|auto_generated|dffe2~q ),
	.dffe17(\u24|u0|auto_generated|dffe1~q ),
	.dffe162(\u24|u0|auto_generated|dffe16~_wirecell_combout ),
	.dffe163(\u27|u0|auto_generated|dffe16~_wirecell_combout ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_cordic_axor_1p_lpm_5 u26(
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.pipeline_dffe_17(\u26|u0|auto_generated|pipeline_dffe[17]~q ),
	.pipeline_dffe_16(\u26|u0|auto_generated|pipeline_dffe[16]~q ),
	.dffe16(\u24|u0|auto_generated|dffe16~q ),
	.pipeline_dffe_15(\u26|u0|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_171(\u23|u0|auto_generated|pipeline_dffe[17]~q ),
	.dffe18(\u22|u0|auto_generated|dffe18~q ),
	.pipeline_dffe_14(\u26|u0|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_13(\u26|u0|auto_generated|pipeline_dffe[13]~q ),
	.dffe17(\u22|u0|auto_generated|dffe17~q ),
	.pipeline_dffe_161(\u23|u0|auto_generated|pipeline_dffe[16]~q ),
	.pipeline_dffe_12(\u26|u0|auto_generated|pipeline_dffe[12]~q ),
	.dffe161(\u22|u0|auto_generated|dffe16~q ),
	.pipeline_dffe_151(\u23|u0|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_11(\u26|u0|auto_generated|pipeline_dffe[11]~q ),
	.dffe15(\u22|u0|auto_generated|dffe15~q ),
	.pipeline_dffe_141(\u23|u0|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_10(\u26|u0|auto_generated|pipeline_dffe[10]~q ),
	.dffe14(\u22|u0|auto_generated|dffe14~q ),
	.pipeline_dffe_9(\u26|u0|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_131(\u23|u0|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_0(\u26|u0|auto_generated|pipeline_dffe[0]~q ),
	.dffe13(\u22|u0|auto_generated|dffe13~q ),
	.pipeline_dffe_121(\u23|u0|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_1(\u26|u0|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_2(\u26|u0|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\u26|u0|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\u26|u0|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\u26|u0|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\u26|u0|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\u26|u0|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\u26|u0|auto_generated|pipeline_dffe[8]~q ),
	.dffe12(\u22|u0|auto_generated|dffe12~q ),
	.pipeline_dffe_111(\u23|u0|auto_generated|pipeline_dffe[11]~q ),
	.dffe11(\u22|u0|auto_generated|dffe11~q ),
	.pipeline_dffe_101(\u23|u0|auto_generated|pipeline_dffe[10]~q ),
	.dffe9(\u22|u0|auto_generated|dffe9~q ),
	.dffe10(\u22|u0|auto_generated|dffe10~q ),
	.pipeline_dffe_81(\u23|u0|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_91(\u23|u0|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_01(\u23|u0|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_18(\u23|u0|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_21(\u23|u0|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_31(\u23|u0|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_41(\u23|u0|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_51(\u23|u0|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_61(\u23|u0|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_71(\u23|u0|auto_generated|pipeline_dffe[7]~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_cordic_sxor_1p_lpm_6 u28(
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.dffe18(\u28|u0|auto_generated|dffe18~q ),
	.dffe17(\u28|u0|auto_generated|dffe17~q ),
	.dffe16(\u27|u0|auto_generated|dffe16~q ),
	.dffe161(\u28|u0|auto_generated|dffe16~q ),
	.dffe181(\u25|u0|auto_generated|dffe18~q ),
	.pipeline_dffe_17(\u26|u0|auto_generated|pipeline_dffe[17]~q ),
	.dffe15(\u28|u0|auto_generated|dffe15~q ),
	.dffe14(\u28|u0|auto_generated|dffe14~q ),
	.pipeline_dffe_16(\u26|u0|auto_generated|pipeline_dffe[16]~q ),
	.dffe171(\u25|u0|auto_generated|dffe17~q ),
	.dffe13(\u28|u0|auto_generated|dffe13~q ),
	.pipeline_dffe_15(\u26|u0|auto_generated|pipeline_dffe[15]~q ),
	.dffe162(\u25|u0|auto_generated|dffe16~q ),
	.dffe11(\u28|u0|auto_generated|dffe11~q ),
	.dffe12(\u28|u0|auto_generated|dffe12~q ),
	.pipeline_dffe_14(\u26|u0|auto_generated|pipeline_dffe[14]~q ),
	.dffe151(\u25|u0|auto_generated|dffe15~q ),
	.pipeline_dffe_13(\u26|u0|auto_generated|pipeline_dffe[13]~q ),
	.dffe1(\u28|u0|auto_generated|dffe1~q ),
	.dffe141(\u25|u0|auto_generated|dffe14~q ),
	.dffe2(\u28|u0|auto_generated|dffe2~q ),
	.dffe3(\u28|u0|auto_generated|dffe3~q ),
	.dffe4(\u28|u0|auto_generated|dffe4~q ),
	.dffe5(\u28|u0|auto_generated|dffe5~q ),
	.dffe6(\u28|u0|auto_generated|dffe6~q ),
	.dffe7(\u28|u0|auto_generated|dffe7~q ),
	.dffe8(\u28|u0|auto_generated|dffe8~q ),
	.dffe9(\u28|u0|auto_generated|dffe9~q ),
	.dffe10(\u28|u0|auto_generated|dffe10~q ),
	.pipeline_dffe_12(\u26|u0|auto_generated|pipeline_dffe[12]~q ),
	.dffe131(\u25|u0|auto_generated|dffe13~q ),
	.pipeline_dffe_11(\u26|u0|auto_generated|pipeline_dffe[11]~q ),
	.dffe121(\u25|u0|auto_generated|dffe12~q ),
	.dffe101(\u25|u0|auto_generated|dffe10~q ),
	.dffe111(\u25|u0|auto_generated|dffe11~q ),
	.pipeline_dffe_10(\u26|u0|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_9(\u26|u0|auto_generated|pipeline_dffe[9]~q ),
	.dffe19(\u25|u0|auto_generated|dffe1~q ),
	.dffe21(\u25|u0|auto_generated|dffe2~q ),
	.dffe31(\u25|u0|auto_generated|dffe3~q ),
	.dffe41(\u25|u0|auto_generated|dffe4~q ),
	.dffe51(\u25|u0|auto_generated|dffe5~q ),
	.dffe61(\u25|u0|auto_generated|dffe6~q ),
	.dffe71(\u25|u0|auto_generated|dffe7~q ),
	.dffe81(\u25|u0|auto_generated|dffe8~q ),
	.dffe91(\u25|u0|auto_generated|dffe9~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_cordic_zxor_1p_lpm_7 u30(
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.dffe16(\u30|u0|auto_generated|dffe16~q ),
	.dffe15(\u30|u0|auto_generated|dffe15~q ),
	.dffe14(\u30|u0|auto_generated|dffe14~q ),
	.dffe161(\u27|u0|auto_generated|dffe16~q ),
	.dffe13(\u30|u0|auto_generated|dffe13~q ),
	.dffe12(\u30|u0|auto_generated|dffe12~q ),
	.dffe151(\u27|u0|auto_generated|dffe15~q ),
	.dffe11(\u30|u0|auto_generated|dffe11~q ),
	.dffe141(\u27|u0|auto_generated|dffe14~q ),
	.dffe10(\u30|u0|auto_generated|dffe10~q ),
	.dffe131(\u27|u0|auto_generated|dffe13~q ),
	.dffe9(\u30|u0|auto_generated|dffe9~q ),
	.dffe121(\u27|u0|auto_generated|dffe12~q ),
	.dffe8(\u30|u0|auto_generated|dffe8~q ),
	.dffe111(\u27|u0|auto_generated|dffe11~q ),
	.dffe7(\u30|u0|auto_generated|dffe7~q ),
	.dffe101(\u27|u0|auto_generated|dffe10~q ),
	.dffe6(\u30|u0|auto_generated|dffe6~q ),
	.dffe91(\u27|u0|auto_generated|dffe9~q ),
	.dffe5(\u30|u0|auto_generated|dffe5~q ),
	.dffe81(\u27|u0|auto_generated|dffe8~q ),
	.dffe4(\u30|u0|auto_generated|dffe4~q ),
	.dffe71(\u27|u0|auto_generated|dffe7~q ),
	.dffe3(\u30|u0|auto_generated|dffe3~q ),
	.dffe61(\u27|u0|auto_generated|dffe6~q ),
	.dffe2(\u30|u0|auto_generated|dffe2~q ),
	.dffe51(\u27|u0|auto_generated|dffe5~q ),
	.dffe1(\u30|u0|auto_generated|dffe1~q ),
	.dffe41(\u27|u0|auto_generated|dffe4~q ),
	.dffe31(\u27|u0|auto_generated|dffe3~q ),
	.dffe21(\u27|u0|auto_generated|dffe2~q ),
	.dffe17(\u27|u0|auto_generated|dffe1~q ),
	.dffe162(\u27|u0|auto_generated|dffe16~_wirecell_combout ),
	.dffe163(\u30|u0|auto_generated|dffe16~_wirecell_combout ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_cordic_axor_1p_lpm_6 u29(
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.pipeline_dffe_17(\u29|u0|auto_generated|pipeline_dffe[17]~q ),
	.pipeline_dffe_16(\u29|u0|auto_generated|pipeline_dffe[16]~q ),
	.dffe16(\u27|u0|auto_generated|dffe16~q ),
	.dffe18(\u25|u0|auto_generated|dffe18~q ),
	.pipeline_dffe_15(\u29|u0|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_171(\u26|u0|auto_generated|pipeline_dffe[17]~q ),
	.pipeline_dffe_14(\u29|u0|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_161(\u26|u0|auto_generated|pipeline_dffe[16]~q ),
	.pipeline_dffe_13(\u29|u0|auto_generated|pipeline_dffe[13]~q ),
	.dffe17(\u25|u0|auto_generated|dffe17~q ),
	.pipeline_dffe_151(\u26|u0|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_12(\u29|u0|auto_generated|pipeline_dffe[12]~q ),
	.dffe161(\u25|u0|auto_generated|dffe16~q ),
	.pipeline_dffe_141(\u26|u0|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_10(\u29|u0|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_11(\u29|u0|auto_generated|pipeline_dffe[11]~q ),
	.dffe15(\u25|u0|auto_generated|dffe15~q ),
	.pipeline_dffe_0(\u29|u0|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_131(\u26|u0|auto_generated|pipeline_dffe[13]~q ),
	.dffe14(\u25|u0|auto_generated|dffe14~q ),
	.pipeline_dffe_1(\u29|u0|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_2(\u29|u0|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\u29|u0|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\u29|u0|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\u29|u0|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\u29|u0|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\u29|u0|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\u29|u0|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\u29|u0|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_121(\u26|u0|auto_generated|pipeline_dffe[12]~q ),
	.dffe13(\u25|u0|auto_generated|dffe13~q ),
	.pipeline_dffe_111(\u26|u0|auto_generated|pipeline_dffe[11]~q ),
	.dffe12(\u25|u0|auto_generated|dffe12~q ),
	.dffe10(\u25|u0|auto_generated|dffe10~q ),
	.dffe11(\u25|u0|auto_generated|dffe11~q ),
	.pipeline_dffe_101(\u26|u0|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_91(\u26|u0|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_01(\u26|u0|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_18(\u26|u0|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_21(\u26|u0|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_31(\u26|u0|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_41(\u26|u0|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_51(\u26|u0|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_61(\u26|u0|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_71(\u26|u0|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_81(\u26|u0|auto_generated|pipeline_dffe[8]~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_cordic_axor_1p_lpm_7 u32(
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.pipeline_dffe_17(\u32|u0|auto_generated|pipeline_dffe[17]~q ),
	.pipeline_dffe_16(\u32|u0|auto_generated|pipeline_dffe[16]~q ),
	.dffe16(\u30|u0|auto_generated|dffe16~q ),
	.pipeline_dffe_15(\u32|u0|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_171(\u29|u0|auto_generated|pipeline_dffe[17]~q ),
	.dffe18(\u28|u0|auto_generated|dffe18~q ),
	.pipeline_dffe_14(\u32|u0|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_13(\u32|u0|auto_generated|pipeline_dffe[13]~q ),
	.dffe17(\u28|u0|auto_generated|dffe17~q ),
	.pipeline_dffe_161(\u29|u0|auto_generated|pipeline_dffe[16]~q ),
	.pipeline_dffe_12(\u32|u0|auto_generated|pipeline_dffe[12]~q ),
	.dffe161(\u28|u0|auto_generated|dffe16~q ),
	.pipeline_dffe_11(\u32|u0|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_151(\u29|u0|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_0(\u32|u0|auto_generated|pipeline_dffe[0]~q ),
	.dffe15(\u28|u0|auto_generated|dffe15~q ),
	.pipeline_dffe_141(\u29|u0|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_1(\u32|u0|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_2(\u32|u0|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\u32|u0|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\u32|u0|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\u32|u0|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\u32|u0|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\u32|u0|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\u32|u0|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\u32|u0|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_10(\u32|u0|auto_generated|pipeline_dffe[10]~q ),
	.dffe14(\u28|u0|auto_generated|dffe14~q ),
	.pipeline_dffe_131(\u29|u0|auto_generated|pipeline_dffe[13]~q ),
	.dffe13(\u28|u0|auto_generated|dffe13~q ),
	.pipeline_dffe_121(\u29|u0|auto_generated|pipeline_dffe[12]~q ),
	.dffe11(\u28|u0|auto_generated|dffe11~q ),
	.dffe12(\u28|u0|auto_generated|dffe12~q ),
	.pipeline_dffe_101(\u29|u0|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_111(\u29|u0|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_01(\u29|u0|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_18(\u29|u0|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_21(\u29|u0|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_31(\u29|u0|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_41(\u29|u0|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_51(\u29|u0|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_61(\u29|u0|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_71(\u29|u0|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_81(\u29|u0|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_91(\u29|u0|auto_generated|pipeline_dffe[9]~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_cordic_sxor_1p_lpm_7 u31(
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.dffe18(\u31|u0|auto_generated|dffe18~q ),
	.dffe17(\u31|u0|auto_generated|dffe17~q ),
	.dffe16(\u30|u0|auto_generated|dffe16~q ),
	.pipeline_dffe_17(\u29|u0|auto_generated|pipeline_dffe[17]~q ),
	.dffe161(\u31|u0|auto_generated|dffe16~q ),
	.dffe181(\u28|u0|auto_generated|dffe18~q ),
	.dffe15(\u31|u0|auto_generated|dffe15~q ),
	.dffe171(\u28|u0|auto_generated|dffe17~q ),
	.dffe14(\u31|u0|auto_generated|dffe14~q ),
	.pipeline_dffe_16(\u29|u0|auto_generated|pipeline_dffe[16]~q ),
	.dffe12(\u31|u0|auto_generated|dffe12~q ),
	.dffe13(\u31|u0|auto_generated|dffe13~q ),
	.dffe162(\u28|u0|auto_generated|dffe16~q ),
	.pipeline_dffe_15(\u29|u0|auto_generated|pipeline_dffe[15]~q ),
	.dffe151(\u28|u0|auto_generated|dffe15~q ),
	.dffe1(\u31|u0|auto_generated|dffe1~q ),
	.pipeline_dffe_14(\u29|u0|auto_generated|pipeline_dffe[14]~q ),
	.dffe2(\u31|u0|auto_generated|dffe2~q ),
	.dffe3(\u31|u0|auto_generated|dffe3~q ),
	.dffe4(\u31|u0|auto_generated|dffe4~q ),
	.dffe5(\u31|u0|auto_generated|dffe5~q ),
	.dffe6(\u31|u0|auto_generated|dffe6~q ),
	.dffe7(\u31|u0|auto_generated|dffe7~q ),
	.dffe8(\u31|u0|auto_generated|dffe8~q ),
	.dffe9(\u31|u0|auto_generated|dffe9~q ),
	.dffe10(\u31|u0|auto_generated|dffe10~q ),
	.dffe11(\u31|u0|auto_generated|dffe11~q ),
	.dffe141(\u28|u0|auto_generated|dffe14~q ),
	.pipeline_dffe_13(\u29|u0|auto_generated|pipeline_dffe[13]~q ),
	.dffe131(\u28|u0|auto_generated|dffe13~q ),
	.pipeline_dffe_12(\u29|u0|auto_generated|pipeline_dffe[12]~q ),
	.dffe111(\u28|u0|auto_generated|dffe11~q ),
	.dffe121(\u28|u0|auto_generated|dffe12~q ),
	.pipeline_dffe_10(\u29|u0|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_11(\u29|u0|auto_generated|pipeline_dffe[11]~q ),
	.dffe19(\u28|u0|auto_generated|dffe1~q ),
	.dffe21(\u28|u0|auto_generated|dffe2~q ),
	.dffe31(\u28|u0|auto_generated|dffe3~q ),
	.dffe41(\u28|u0|auto_generated|dffe4~q ),
	.dffe51(\u28|u0|auto_generated|dffe5~q ),
	.dffe61(\u28|u0|auto_generated|dffe6~q ),
	.dffe71(\u28|u0|auto_generated|dffe7~q ),
	.dffe81(\u28|u0|auto_generated|dffe8~q ),
	.dffe91(\u28|u0|auto_generated|dffe9~q ),
	.dffe101(\u28|u0|auto_generated|dffe10~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_cordic_sxor_1p_lpm_8 u34(
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.dffe18(\u34|u0|auto_generated|dffe18~q ),
	.dffe17(\u34|u0|auto_generated|dffe17~q ),
	.dffe16(\u33|u0|auto_generated|dffe16~q ),
	.dffe161(\u34|u0|auto_generated|dffe16~q ),
	.dffe181(\u31|u0|auto_generated|dffe18~q ),
	.pipeline_dffe_17(\u32|u0|auto_generated|pipeline_dffe[17]~q ),
	.dffe15(\u34|u0|auto_generated|dffe15~q ),
	.dffe13(\u34|u0|auto_generated|dffe13~q ),
	.dffe14(\u34|u0|auto_generated|dffe14~q ),
	.pipeline_dffe_16(\u32|u0|auto_generated|pipeline_dffe[16]~q ),
	.dffe171(\u31|u0|auto_generated|dffe17~q ),
	.pipeline_dffe_15(\u32|u0|auto_generated|pipeline_dffe[15]~q ),
	.dffe1(\u34|u0|auto_generated|dffe1~q ),
	.dffe162(\u31|u0|auto_generated|dffe16~q ),
	.dffe2(\u34|u0|auto_generated|dffe2~q ),
	.dffe3(\u34|u0|auto_generated|dffe3~q ),
	.dffe4(\u34|u0|auto_generated|dffe4~q ),
	.dffe5(\u34|u0|auto_generated|dffe5~q ),
	.dffe6(\u34|u0|auto_generated|dffe6~q ),
	.dffe7(\u34|u0|auto_generated|dffe7~q ),
	.dffe8(\u34|u0|auto_generated|dffe8~q ),
	.dffe9(\u34|u0|auto_generated|dffe9~q ),
	.dffe10(\u34|u0|auto_generated|dffe10~q ),
	.dffe11(\u34|u0|auto_generated|dffe11~q ),
	.dffe12(\u34|u0|auto_generated|dffe12~q ),
	.pipeline_dffe_14(\u32|u0|auto_generated|pipeline_dffe[14]~q ),
	.dffe151(\u31|u0|auto_generated|dffe15~q ),
	.pipeline_dffe_13(\u32|u0|auto_generated|pipeline_dffe[13]~q ),
	.dffe141(\u31|u0|auto_generated|dffe14~q ),
	.dffe121(\u31|u0|auto_generated|dffe12~q ),
	.dffe131(\u31|u0|auto_generated|dffe13~q ),
	.pipeline_dffe_12(\u32|u0|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_11(\u32|u0|auto_generated|pipeline_dffe[11]~q ),
	.dffe19(\u31|u0|auto_generated|dffe1~q ),
	.dffe21(\u31|u0|auto_generated|dffe2~q ),
	.dffe31(\u31|u0|auto_generated|dffe3~q ),
	.dffe41(\u31|u0|auto_generated|dffe4~q ),
	.dffe51(\u31|u0|auto_generated|dffe5~q ),
	.dffe61(\u31|u0|auto_generated|dffe6~q ),
	.dffe71(\u31|u0|auto_generated|dffe7~q ),
	.dffe81(\u31|u0|auto_generated|dffe8~q ),
	.dffe91(\u31|u0|auto_generated|dffe9~q ),
	.dffe101(\u31|u0|auto_generated|dffe10~q ),
	.dffe111(\u31|u0|auto_generated|dffe11~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_cordic_zxor_1p_lpm_8 u33(
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.dffe16(\u33|u0|auto_generated|dffe16~q ),
	.dffe15(\u33|u0|auto_generated|dffe15~q ),
	.dffe14(\u33|u0|auto_generated|dffe14~q ),
	.dffe161(\u30|u0|auto_generated|dffe16~q ),
	.dffe13(\u33|u0|auto_generated|dffe13~q ),
	.dffe12(\u33|u0|auto_generated|dffe12~q ),
	.dffe151(\u30|u0|auto_generated|dffe15~q ),
	.dffe11(\u33|u0|auto_generated|dffe11~q ),
	.dffe141(\u30|u0|auto_generated|dffe14~q ),
	.dffe10(\u33|u0|auto_generated|dffe10~q ),
	.dffe131(\u30|u0|auto_generated|dffe13~q ),
	.dffe9(\u33|u0|auto_generated|dffe9~q ),
	.dffe121(\u30|u0|auto_generated|dffe12~q ),
	.dffe8(\u33|u0|auto_generated|dffe8~q ),
	.dffe111(\u30|u0|auto_generated|dffe11~q ),
	.dffe7(\u33|u0|auto_generated|dffe7~q ),
	.dffe101(\u30|u0|auto_generated|dffe10~q ),
	.dffe6(\u33|u0|auto_generated|dffe6~q ),
	.dffe91(\u30|u0|auto_generated|dffe9~q ),
	.dffe5(\u33|u0|auto_generated|dffe5~q ),
	.dffe81(\u30|u0|auto_generated|dffe8~q ),
	.dffe4(\u33|u0|auto_generated|dffe4~q ),
	.dffe71(\u30|u0|auto_generated|dffe7~q ),
	.dffe3(\u33|u0|auto_generated|dffe3~q ),
	.dffe61(\u30|u0|auto_generated|dffe6~q ),
	.dffe2(\u33|u0|auto_generated|dffe2~q ),
	.dffe51(\u30|u0|auto_generated|dffe5~q ),
	.dffe1(\u33|u0|auto_generated|dffe1~q ),
	.dffe41(\u30|u0|auto_generated|dffe4~q ),
	.dffe31(\u30|u0|auto_generated|dffe3~q ),
	.dffe21(\u30|u0|auto_generated|dffe2~q ),
	.dffe17(\u30|u0|auto_generated|dffe1~q ),
	.dffe162(\u30|u0|auto_generated|dffe16~_wirecell_combout ),
	.dffe163(\u33|u0|auto_generated|dffe16~_wirecell_combout ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_cordic_zxor_1p_lpm_9 u36(
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.dffe16(\u36|u0|auto_generated|dffe16~q ),
	.dffe15(\u36|u0|auto_generated|dffe15~q ),
	.dffe14(\u36|u0|auto_generated|dffe14~q ),
	.dffe161(\u33|u0|auto_generated|dffe16~q ),
	.dffe13(\u36|u0|auto_generated|dffe13~q ),
	.dffe12(\u36|u0|auto_generated|dffe12~q ),
	.dffe151(\u33|u0|auto_generated|dffe15~q ),
	.dffe11(\u36|u0|auto_generated|dffe11~q ),
	.dffe141(\u33|u0|auto_generated|dffe14~q ),
	.dffe10(\u36|u0|auto_generated|dffe10~q ),
	.dffe131(\u33|u0|auto_generated|dffe13~q ),
	.dffe9(\u36|u0|auto_generated|dffe9~q ),
	.dffe121(\u33|u0|auto_generated|dffe12~q ),
	.dffe8(\u36|u0|auto_generated|dffe8~q ),
	.dffe111(\u33|u0|auto_generated|dffe11~q ),
	.dffe7(\u36|u0|auto_generated|dffe7~q ),
	.dffe101(\u33|u0|auto_generated|dffe10~q ),
	.dffe6(\u36|u0|auto_generated|dffe6~q ),
	.dffe91(\u33|u0|auto_generated|dffe9~q ),
	.dffe5(\u36|u0|auto_generated|dffe5~q ),
	.dffe81(\u33|u0|auto_generated|dffe8~q ),
	.dffe4(\u36|u0|auto_generated|dffe4~q ),
	.dffe71(\u33|u0|auto_generated|dffe7~q ),
	.dffe3(\u36|u0|auto_generated|dffe3~q ),
	.dffe61(\u33|u0|auto_generated|dffe6~q ),
	.dffe2(\u36|u0|auto_generated|dffe2~q ),
	.dffe51(\u33|u0|auto_generated|dffe5~q ),
	.dffe1(\u36|u0|auto_generated|dffe1~q ),
	.dffe41(\u33|u0|auto_generated|dffe4~q ),
	.dffe31(\u33|u0|auto_generated|dffe3~q ),
	.dffe21(\u33|u0|auto_generated|dffe2~q ),
	.dffe17(\u33|u0|auto_generated|dffe1~q ),
	.dffe162(\u33|u0|auto_generated|dffe16~_wirecell_combout ),
	.dffe163(\u36|u0|auto_generated|dffe16~_wirecell_combout ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_cordic_axor_1p_lpm_8 u35(
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.pipeline_dffe_17(\u35|u0|auto_generated|pipeline_dffe[17]~q ),
	.pipeline_dffe_16(\u35|u0|auto_generated|pipeline_dffe[16]~q ),
	.dffe16(\u33|u0|auto_generated|dffe16~q ),
	.dffe18(\u31|u0|auto_generated|dffe18~q ),
	.pipeline_dffe_15(\u35|u0|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_171(\u32|u0|auto_generated|pipeline_dffe[17]~q ),
	.pipeline_dffe_14(\u35|u0|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_161(\u32|u0|auto_generated|pipeline_dffe[16]~q ),
	.pipeline_dffe_12(\u35|u0|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_13(\u35|u0|auto_generated|pipeline_dffe[13]~q ),
	.dffe17(\u31|u0|auto_generated|dffe17~q ),
	.pipeline_dffe_0(\u35|u0|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_151(\u32|u0|auto_generated|pipeline_dffe[15]~q ),
	.dffe161(\u31|u0|auto_generated|dffe16~q ),
	.pipeline_dffe_1(\u35|u0|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_2(\u35|u0|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\u35|u0|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\u35|u0|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\u35|u0|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\u35|u0|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\u35|u0|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\u35|u0|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\u35|u0|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_10(\u35|u0|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_11(\u35|u0|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_141(\u32|u0|auto_generated|pipeline_dffe[14]~q ),
	.dffe15(\u31|u0|auto_generated|dffe15~q ),
	.pipeline_dffe_131(\u32|u0|auto_generated|pipeline_dffe[13]~q ),
	.dffe14(\u31|u0|auto_generated|dffe14~q ),
	.dffe12(\u31|u0|auto_generated|dffe12~q ),
	.dffe13(\u31|u0|auto_generated|dffe13~q ),
	.pipeline_dffe_121(\u32|u0|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_111(\u32|u0|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_01(\u32|u0|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_18(\u32|u0|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_21(\u32|u0|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_31(\u32|u0|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_41(\u32|u0|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_51(\u32|u0|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_61(\u32|u0|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_71(\u32|u0|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_81(\u32|u0|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_91(\u32|u0|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_101(\u32|u0|auto_generated|pipeline_dffe[10]~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_cordic_axor_1p_lpm_9 u38(
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.pipeline_dffe_17(\u38|u0|auto_generated|pipeline_dffe[17]~q ),
	.pipeline_dffe_16(\u38|u0|auto_generated|pipeline_dffe[16]~q ),
	.dffe16(\u36|u0|auto_generated|dffe16~q ),
	.pipeline_dffe_15(\u38|u0|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_171(\u35|u0|auto_generated|pipeline_dffe[17]~q ),
	.dffe18(\u34|u0|auto_generated|dffe18~q ),
	.pipeline_dffe_14(\u38|u0|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_13(\u38|u0|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_0(\u38|u0|auto_generated|pipeline_dffe[0]~q ),
	.dffe17(\u34|u0|auto_generated|dffe17~q ),
	.pipeline_dffe_161(\u35|u0|auto_generated|pipeline_dffe[16]~q ),
	.pipeline_dffe_1(\u38|u0|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_2(\u38|u0|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\u38|u0|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\u38|u0|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\u38|u0|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\u38|u0|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\u38|u0|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\u38|u0|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\u38|u0|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_10(\u38|u0|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_11(\u38|u0|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_12(\u38|u0|auto_generated|pipeline_dffe[12]~q ),
	.dffe161(\u34|u0|auto_generated|dffe16~q ),
	.pipeline_dffe_151(\u35|u0|auto_generated|pipeline_dffe[15]~q ),
	.dffe15(\u34|u0|auto_generated|dffe15~q ),
	.pipeline_dffe_141(\u35|u0|auto_generated|pipeline_dffe[14]~q ),
	.dffe13(\u34|u0|auto_generated|dffe13~q ),
	.dffe14(\u34|u0|auto_generated|dffe14~q ),
	.pipeline_dffe_121(\u35|u0|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_131(\u35|u0|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_01(\u35|u0|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_18(\u35|u0|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_21(\u35|u0|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_31(\u35|u0|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_41(\u35|u0|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_51(\u35|u0|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_61(\u35|u0|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_71(\u35|u0|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_81(\u35|u0|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_91(\u35|u0|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_101(\u35|u0|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_111(\u35|u0|auto_generated|pipeline_dffe[11]~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_cordic_sxor_1p_lpm_9 u37(
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.dffe18(\u37|u0|auto_generated|dffe18~q ),
	.dffe17(\u37|u0|auto_generated|dffe17~q ),
	.dffe16(\u36|u0|auto_generated|dffe16~q ),
	.pipeline_dffe_17(\u35|u0|auto_generated|pipeline_dffe[17]~q ),
	.dffe161(\u37|u0|auto_generated|dffe16~q ),
	.dffe181(\u34|u0|auto_generated|dffe18~q ),
	.dffe14(\u37|u0|auto_generated|dffe14~q ),
	.dffe15(\u37|u0|auto_generated|dffe15~q ),
	.dffe171(\u34|u0|auto_generated|dffe17~q ),
	.dffe1(\u37|u0|auto_generated|dffe1~q ),
	.pipeline_dffe_16(\u35|u0|auto_generated|pipeline_dffe[16]~q ),
	.dffe2(\u37|u0|auto_generated|dffe2~q ),
	.dffe3(\u37|u0|auto_generated|dffe3~q ),
	.dffe4(\u37|u0|auto_generated|dffe4~q ),
	.dffe5(\u37|u0|auto_generated|dffe5~q ),
	.dffe6(\u37|u0|auto_generated|dffe6~q ),
	.dffe7(\u37|u0|auto_generated|dffe7~q ),
	.dffe8(\u37|u0|auto_generated|dffe8~q ),
	.dffe9(\u37|u0|auto_generated|dffe9~q ),
	.dffe10(\u37|u0|auto_generated|dffe10~q ),
	.dffe11(\u37|u0|auto_generated|dffe11~q ),
	.dffe12(\u37|u0|auto_generated|dffe12~q ),
	.dffe13(\u37|u0|auto_generated|dffe13~q ),
	.dffe162(\u34|u0|auto_generated|dffe16~q ),
	.pipeline_dffe_15(\u35|u0|auto_generated|pipeline_dffe[15]~q ),
	.dffe151(\u34|u0|auto_generated|dffe15~q ),
	.pipeline_dffe_14(\u35|u0|auto_generated|pipeline_dffe[14]~q ),
	.dffe131(\u34|u0|auto_generated|dffe13~q ),
	.dffe141(\u34|u0|auto_generated|dffe14~q ),
	.pipeline_dffe_12(\u35|u0|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_13(\u35|u0|auto_generated|pipeline_dffe[13]~q ),
	.dffe19(\u34|u0|auto_generated|dffe1~q ),
	.dffe21(\u34|u0|auto_generated|dffe2~q ),
	.dffe31(\u34|u0|auto_generated|dffe3~q ),
	.dffe41(\u34|u0|auto_generated|dffe4~q ),
	.dffe51(\u34|u0|auto_generated|dffe5~q ),
	.dffe61(\u34|u0|auto_generated|dffe6~q ),
	.dffe71(\u34|u0|auto_generated|dffe7~q ),
	.dffe81(\u34|u0|auto_generated|dffe8~q ),
	.dffe91(\u34|u0|auto_generated|dffe9~q ),
	.dffe101(\u34|u0|auto_generated|dffe10~q ),
	.dffe111(\u34|u0|auto_generated|dffe11~q ),
	.dffe121(\u34|u0|auto_generated|dffe12~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_cordic_sxor_1p_lpm_11 u40(
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.dffe18(\u40|u0|auto_generated|dffe18~q ),
	.dffe17(\u40|u0|auto_generated|dffe17~q ),
	.dffe15(\u40|u0|auto_generated|dffe15~q ),
	.dffe16(\u40|u0|auto_generated|dffe16~q ),
	.dffe161(\u39|u0|auto_generated|dffe16~q ),
	.dffe181(\u37|u0|auto_generated|dffe18~q ),
	.pipeline_dffe_17(\u38|u0|auto_generated|pipeline_dffe[17]~q ),
	.dffe1(\u40|u0|auto_generated|dffe1~q ),
	.dffe2(\u40|u0|auto_generated|dffe2~q ),
	.dffe3(\u40|u0|auto_generated|dffe3~q ),
	.dffe4(\u40|u0|auto_generated|dffe4~q ),
	.dffe5(\u40|u0|auto_generated|dffe5~q ),
	.dffe6(\u40|u0|auto_generated|dffe6~q ),
	.dffe7(\u40|u0|auto_generated|dffe7~q ),
	.dffe8(\u40|u0|auto_generated|dffe8~q ),
	.dffe9(\u40|u0|auto_generated|dffe9~q ),
	.dffe10(\u40|u0|auto_generated|dffe10~q ),
	.dffe11(\u40|u0|auto_generated|dffe11~q ),
	.dffe12(\u40|u0|auto_generated|dffe12~q ),
	.dffe13(\u40|u0|auto_generated|dffe13~q ),
	.dffe14(\u40|u0|auto_generated|dffe14~q ),
	.pipeline_dffe_16(\u38|u0|auto_generated|pipeline_dffe[16]~q ),
	.dffe171(\u37|u0|auto_generated|dffe17~q ),
	.pipeline_dffe_15(\u38|u0|auto_generated|pipeline_dffe[15]~q ),
	.dffe162(\u37|u0|auto_generated|dffe16~q ),
	.dffe141(\u37|u0|auto_generated|dffe14~q ),
	.dffe151(\u37|u0|auto_generated|dffe15~q ),
	.pipeline_dffe_14(\u38|u0|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_13(\u38|u0|auto_generated|pipeline_dffe[13]~q ),
	.dffe19(\u37|u0|auto_generated|dffe1~q ),
	.dffe21(\u37|u0|auto_generated|dffe2~q ),
	.dffe31(\u37|u0|auto_generated|dffe3~q ),
	.dffe41(\u37|u0|auto_generated|dffe4~q ),
	.dffe51(\u37|u0|auto_generated|dffe5~q ),
	.dffe61(\u37|u0|auto_generated|dffe6~q ),
	.dffe71(\u37|u0|auto_generated|dffe7~q ),
	.dffe81(\u37|u0|auto_generated|dffe8~q ),
	.dffe91(\u37|u0|auto_generated|dffe9~q ),
	.dffe101(\u37|u0|auto_generated|dffe10~q ),
	.dffe111(\u37|u0|auto_generated|dffe11~q ),
	.dffe121(\u37|u0|auto_generated|dffe12~q ),
	.dffe131(\u37|u0|auto_generated|dffe13~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_cordic_zxor_1p_lpm_10 u39(
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.dffe16(\u39|u0|auto_generated|dffe16~q ),
	.dffe15(\u39|u0|auto_generated|dffe15~q ),
	.dffe14(\u39|u0|auto_generated|dffe14~q ),
	.dffe161(\u36|u0|auto_generated|dffe16~q ),
	.dffe13(\u39|u0|auto_generated|dffe13~q ),
	.dffe12(\u39|u0|auto_generated|dffe12~q ),
	.dffe151(\u36|u0|auto_generated|dffe15~q ),
	.dffe11(\u39|u0|auto_generated|dffe11~q ),
	.dffe141(\u36|u0|auto_generated|dffe14~q ),
	.dffe10(\u39|u0|auto_generated|dffe10~q ),
	.dffe131(\u36|u0|auto_generated|dffe13~q ),
	.dffe9(\u39|u0|auto_generated|dffe9~q ),
	.dffe121(\u36|u0|auto_generated|dffe12~q ),
	.dffe8(\u39|u0|auto_generated|dffe8~q ),
	.dffe111(\u36|u0|auto_generated|dffe11~q ),
	.dffe7(\u39|u0|auto_generated|dffe7~q ),
	.dffe101(\u36|u0|auto_generated|dffe10~q ),
	.dffe6(\u39|u0|auto_generated|dffe6~q ),
	.dffe91(\u36|u0|auto_generated|dffe9~q ),
	.dffe5(\u39|u0|auto_generated|dffe5~q ),
	.dffe81(\u36|u0|auto_generated|dffe8~q ),
	.dffe4(\u39|u0|auto_generated|dffe4~q ),
	.dffe71(\u36|u0|auto_generated|dffe7~q ),
	.dffe3(\u39|u0|auto_generated|dffe3~q ),
	.dffe61(\u36|u0|auto_generated|dffe6~q ),
	.dffe2(\u39|u0|auto_generated|dffe2~q ),
	.dffe51(\u36|u0|auto_generated|dffe5~q ),
	.dffe1(\u39|u0|auto_generated|dffe1~q ),
	.dffe41(\u36|u0|auto_generated|dffe4~q ),
	.dffe31(\u36|u0|auto_generated|dffe3~q ),
	.dffe21(\u36|u0|auto_generated|dffe2~q ),
	.dffe17(\u36|u0|auto_generated|dffe1~q ),
	.dffe162(\u36|u0|auto_generated|dffe16~_wirecell_combout ),
	.dffe163(\u39|u0|auto_generated|dffe16~_wirecell_combout ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_cordic_zxor_1p_lpm_11 u42(
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.dffe16(\u42|u0|auto_generated|dffe16~q ),
	.dffe15(\u42|u0|auto_generated|dffe15~q ),
	.dffe14(\u42|u0|auto_generated|dffe14~q ),
	.dffe161(\u39|u0|auto_generated|dffe16~q ),
	.dffe13(\u42|u0|auto_generated|dffe13~q ),
	.dffe12(\u42|u0|auto_generated|dffe12~q ),
	.dffe151(\u39|u0|auto_generated|dffe15~q ),
	.dffe11(\u42|u0|auto_generated|dffe11~q ),
	.dffe141(\u39|u0|auto_generated|dffe14~q ),
	.dffe10(\u42|u0|auto_generated|dffe10~q ),
	.dffe131(\u39|u0|auto_generated|dffe13~q ),
	.dffe9(\u42|u0|auto_generated|dffe9~q ),
	.dffe121(\u39|u0|auto_generated|dffe12~q ),
	.dffe8(\u42|u0|auto_generated|dffe8~q ),
	.dffe111(\u39|u0|auto_generated|dffe11~q ),
	.dffe7(\u42|u0|auto_generated|dffe7~q ),
	.dffe101(\u39|u0|auto_generated|dffe10~q ),
	.dffe6(\u42|u0|auto_generated|dffe6~q ),
	.dffe91(\u39|u0|auto_generated|dffe9~q ),
	.dffe5(\u42|u0|auto_generated|dffe5~q ),
	.dffe81(\u39|u0|auto_generated|dffe8~q ),
	.dffe4(\u42|u0|auto_generated|dffe4~q ),
	.dffe71(\u39|u0|auto_generated|dffe7~q ),
	.dffe3(\u42|u0|auto_generated|dffe3~q ),
	.dffe61(\u39|u0|auto_generated|dffe6~q ),
	.dffe2(\u42|u0|auto_generated|dffe2~q ),
	.dffe51(\u39|u0|auto_generated|dffe5~q ),
	.dffe1(\u42|u0|auto_generated|dffe1~q ),
	.dffe41(\u39|u0|auto_generated|dffe4~q ),
	.dffe31(\u39|u0|auto_generated|dffe3~q ),
	.dffe21(\u39|u0|auto_generated|dffe2~q ),
	.dffe17(\u39|u0|auto_generated|dffe1~q ),
	.dffe162(\u39|u0|auto_generated|dffe16~_wirecell_combout ),
	.dffe163(\u42|u0|auto_generated|dffe16~_wirecell_combout ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_cordic_axor_1p_lpm_10 u41(
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.pipeline_dffe_17(\u41|u0|auto_generated|pipeline_dffe[17]~q ),
	.pipeline_dffe_16(\u41|u0|auto_generated|pipeline_dffe[16]~q ),
	.dffe16(\u39|u0|auto_generated|dffe16~q ),
	.dffe18(\u37|u0|auto_generated|dffe18~q ),
	.pipeline_dffe_14(\u41|u0|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_15(\u41|u0|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_171(\u38|u0|auto_generated|pipeline_dffe[17]~q ),
	.pipeline_dffe_0(\u41|u0|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_1(\u41|u0|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_2(\u41|u0|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\u41|u0|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\u41|u0|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\u41|u0|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\u41|u0|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\u41|u0|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\u41|u0|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\u41|u0|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_10(\u41|u0|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_11(\u41|u0|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_12(\u41|u0|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_13(\u41|u0|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_161(\u38|u0|auto_generated|pipeline_dffe[16]~q ),
	.dffe17(\u37|u0|auto_generated|dffe17~q ),
	.pipeline_dffe_151(\u38|u0|auto_generated|pipeline_dffe[15]~q ),
	.dffe161(\u37|u0|auto_generated|dffe16~q ),
	.dffe14(\u37|u0|auto_generated|dffe14~q ),
	.dffe15(\u37|u0|auto_generated|dffe15~q ),
	.pipeline_dffe_141(\u38|u0|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_131(\u38|u0|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_01(\u38|u0|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_18(\u38|u0|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_21(\u38|u0|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_31(\u38|u0|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_41(\u38|u0|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_51(\u38|u0|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_61(\u38|u0|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_71(\u38|u0|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_81(\u38|u0|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_91(\u38|u0|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_101(\u38|u0|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_111(\u38|u0|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_121(\u38|u0|auto_generated|pipeline_dffe[12]~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_cordic_sxor_1p_lpm_12 u43(
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.dffe18(\u43|u0|auto_generated|dffe18~q ),
	.dffe16(\u43|u0|auto_generated|dffe16~q ),
	.dffe17(\u43|u0|auto_generated|dffe17~q ),
	.dffe161(\u42|u0|auto_generated|dffe16~q ),
	.pipeline_dffe_17(\u41|u0|auto_generated|pipeline_dffe[17]~q ),
	.dffe1(\u43|u0|auto_generated|dffe1~q ),
	.dffe181(\u40|u0|auto_generated|dffe18~q ),
	.dffe2(\u43|u0|auto_generated|dffe2~q ),
	.dffe3(\u43|u0|auto_generated|dffe3~q ),
	.dffe4(\u43|u0|auto_generated|dffe4~q ),
	.dffe5(\u43|u0|auto_generated|dffe5~q ),
	.dffe6(\u43|u0|auto_generated|dffe6~q ),
	.dffe7(\u43|u0|auto_generated|dffe7~q ),
	.dffe8(\u43|u0|auto_generated|dffe8~q ),
	.dffe9(\u43|u0|auto_generated|dffe9~q ),
	.dffe10(\u43|u0|auto_generated|dffe10~q ),
	.dffe11(\u43|u0|auto_generated|dffe11~q ),
	.dffe12(\u43|u0|auto_generated|dffe12~q ),
	.dffe13(\u43|u0|auto_generated|dffe13~q ),
	.dffe14(\u43|u0|auto_generated|dffe14~q ),
	.dffe15(\u43|u0|auto_generated|dffe15~q ),
	.dffe171(\u40|u0|auto_generated|dffe17~q ),
	.pipeline_dffe_16(\u41|u0|auto_generated|pipeline_dffe[16]~q ),
	.dffe151(\u40|u0|auto_generated|dffe15~q ),
	.dffe162(\u40|u0|auto_generated|dffe16~q ),
	.pipeline_dffe_14(\u41|u0|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_15(\u41|u0|auto_generated|pipeline_dffe[15]~q ),
	.dffe19(\u40|u0|auto_generated|dffe1~q ),
	.dffe21(\u40|u0|auto_generated|dffe2~q ),
	.dffe31(\u40|u0|auto_generated|dffe3~q ),
	.dffe41(\u40|u0|auto_generated|dffe4~q ),
	.dffe51(\u40|u0|auto_generated|dffe5~q ),
	.dffe61(\u40|u0|auto_generated|dffe6~q ),
	.dffe71(\u40|u0|auto_generated|dffe7~q ),
	.dffe81(\u40|u0|auto_generated|dffe8~q ),
	.dffe91(\u40|u0|auto_generated|dffe9~q ),
	.dffe101(\u40|u0|auto_generated|dffe10~q ),
	.dffe111(\u40|u0|auto_generated|dffe11~q ),
	.dffe121(\u40|u0|auto_generated|dffe12~q ),
	.dffe131(\u40|u0|auto_generated|dffe13~q ),
	.dffe141(\u40|u0|auto_generated|dffe14~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_cordic_zxor_1p_lpm_12 u45(
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.dffe16(\u45|u0|auto_generated|dffe16~q ),
	.dffe15(\u45|u0|auto_generated|dffe15~q ),
	.dffe14(\u45|u0|auto_generated|dffe14~q ),
	.dffe161(\u42|u0|auto_generated|dffe16~q ),
	.dffe13(\u45|u0|auto_generated|dffe13~q ),
	.dffe12(\u45|u0|auto_generated|dffe12~q ),
	.dffe151(\u42|u0|auto_generated|dffe15~q ),
	.dffe11(\u45|u0|auto_generated|dffe11~q ),
	.dffe141(\u42|u0|auto_generated|dffe14~q ),
	.dffe10(\u45|u0|auto_generated|dffe10~q ),
	.dffe131(\u42|u0|auto_generated|dffe13~q ),
	.dffe9(\u45|u0|auto_generated|dffe9~q ),
	.dffe121(\u42|u0|auto_generated|dffe12~q ),
	.dffe8(\u45|u0|auto_generated|dffe8~q ),
	.dffe111(\u42|u0|auto_generated|dffe11~q ),
	.dffe7(\u45|u0|auto_generated|dffe7~q ),
	.dffe101(\u42|u0|auto_generated|dffe10~q ),
	.dffe6(\u45|u0|auto_generated|dffe6~q ),
	.dffe91(\u42|u0|auto_generated|dffe9~q ),
	.dffe5(\u45|u0|auto_generated|dffe5~q ),
	.dffe81(\u42|u0|auto_generated|dffe8~q ),
	.dffe4(\u45|u0|auto_generated|dffe4~q ),
	.dffe71(\u42|u0|auto_generated|dffe7~q ),
	.dffe3(\u45|u0|auto_generated|dffe3~q ),
	.dffe61(\u42|u0|auto_generated|dffe6~q ),
	.dffe2(\u45|u0|auto_generated|dffe2~q ),
	.dffe51(\u42|u0|auto_generated|dffe5~q ),
	.dffe1(\u45|u0|auto_generated|dffe1~q ),
	.dffe41(\u42|u0|auto_generated|dffe4~q ),
	.dffe31(\u42|u0|auto_generated|dffe3~q ),
	.dffe21(\u42|u0|auto_generated|dffe2~q ),
	.dffe17(\u42|u0|auto_generated|dffe1~q ),
	.dffe162(\u42|u0|auto_generated|dffe16~_wirecell_combout ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_cordic_axor_1p_lpm_11 u44(
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.pipeline_dffe_17(\u44|u0|auto_generated|pipeline_dffe[17]~q ),
	.pipeline_dffe_16(\u44|u0|auto_generated|pipeline_dffe[16]~q ),
	.pipeline_dffe_15(\u44|u0|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_0(\u44|u0|auto_generated|pipeline_dffe[0]~q ),
	.dffe16(\u42|u0|auto_generated|dffe16~q ),
	.pipeline_dffe_171(\u41|u0|auto_generated|pipeline_dffe[17]~q ),
	.dffe18(\u40|u0|auto_generated|dffe18~q ),
	.pipeline_dffe_1(\u44|u0|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_2(\u44|u0|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\u44|u0|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\u44|u0|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\u44|u0|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\u44|u0|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\u44|u0|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\u44|u0|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\u44|u0|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_10(\u44|u0|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_11(\u44|u0|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_12(\u44|u0|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_13(\u44|u0|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_14(\u44|u0|auto_generated|pipeline_dffe[14]~q ),
	.dffe17(\u40|u0|auto_generated|dffe17~q ),
	.pipeline_dffe_161(\u41|u0|auto_generated|pipeline_dffe[16]~q ),
	.dffe15(\u40|u0|auto_generated|dffe15~q ),
	.dffe161(\u40|u0|auto_generated|dffe16~q ),
	.pipeline_dffe_141(\u41|u0|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_151(\u41|u0|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_01(\u41|u0|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_18(\u41|u0|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_21(\u41|u0|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_31(\u41|u0|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_41(\u41|u0|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_51(\u41|u0|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_61(\u41|u0|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_71(\u41|u0|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_81(\u41|u0|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_91(\u41|u0|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_101(\u41|u0|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_111(\u41|u0|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_121(\u41|u0|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_131(\u41|u0|auto_generated|pipeline_dffe[13]~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_cordic_axor_1p_lpm_12 u47(
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.pipeline_dffe_17(\u47|u0|auto_generated|pipeline_dffe[17]~q ),
	.pipeline_dffe_16(\u47|u0|auto_generated|pipeline_dffe[16]~q ),
	.pipeline_dffe_0(\u47|u0|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_1(\u47|u0|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_2(\u47|u0|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\u47|u0|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\u47|u0|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\u47|u0|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\u47|u0|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\u47|u0|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\u47|u0|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\u47|u0|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_10(\u47|u0|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_11(\u47|u0|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_12(\u47|u0|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_13(\u47|u0|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_14(\u47|u0|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_15(\u47|u0|auto_generated|pipeline_dffe[15]~q ),
	.dffe16(\u45|u0|auto_generated|dffe16~q ),
	.dffe18(\u43|u0|auto_generated|dffe18~q ),
	.pipeline_dffe_171(\u44|u0|auto_generated|pipeline_dffe[17]~q ),
	.dffe161(\u43|u0|auto_generated|dffe16~q ),
	.dffe17(\u43|u0|auto_generated|dffe17~q ),
	.pipeline_dffe_161(\u44|u0|auto_generated|pipeline_dffe[16]~q ),
	.pipeline_dffe_151(\u44|u0|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_01(\u44|u0|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_18(\u44|u0|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_21(\u44|u0|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_31(\u44|u0|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_41(\u44|u0|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_51(\u44|u0|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_61(\u44|u0|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_71(\u44|u0|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_81(\u44|u0|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_91(\u44|u0|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_101(\u44|u0|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_111(\u44|u0|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_121(\u44|u0|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_131(\u44|u0|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_141(\u44|u0|auto_generated|pipeline_dffe[14]~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_cordic_sxor_1p_lpm_13 u46(
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.dffe18(\u46|u0|auto_generated|dffe18~q ),
	.dffe17(\u46|u0|auto_generated|dffe17~q ),
	.dffe1(\u46|u0|auto_generated|dffe1~q ),
	.dffe2(\u46|u0|auto_generated|dffe2~q ),
	.dffe3(\u46|u0|auto_generated|dffe3~q ),
	.dffe4(\u46|u0|auto_generated|dffe4~q ),
	.dffe5(\u46|u0|auto_generated|dffe5~q ),
	.dffe6(\u46|u0|auto_generated|dffe6~q ),
	.dffe7(\u46|u0|auto_generated|dffe7~q ),
	.dffe8(\u46|u0|auto_generated|dffe8~q ),
	.dffe9(\u46|u0|auto_generated|dffe9~q ),
	.dffe10(\u46|u0|auto_generated|dffe10~q ),
	.dffe11(\u46|u0|auto_generated|dffe11~q ),
	.dffe12(\u46|u0|auto_generated|dffe12~q ),
	.dffe13(\u46|u0|auto_generated|dffe13~q ),
	.dffe14(\u46|u0|auto_generated|dffe14~q ),
	.dffe15(\u46|u0|auto_generated|dffe15~q ),
	.dffe16(\u46|u0|auto_generated|dffe16~q ),
	.dffe161(\u45|u0|auto_generated|dffe16~q ),
	.dffe181(\u43|u0|auto_generated|dffe18~q ),
	.pipeline_dffe_17(\u44|u0|auto_generated|pipeline_dffe[17]~q ),
	.dffe162(\u43|u0|auto_generated|dffe16~q ),
	.dffe171(\u43|u0|auto_generated|dffe17~q ),
	.pipeline_dffe_16(\u44|u0|auto_generated|pipeline_dffe[16]~q ),
	.pipeline_dffe_15(\u44|u0|auto_generated|pipeline_dffe[15]~q ),
	.dffe19(\u43|u0|auto_generated|dffe1~q ),
	.dffe21(\u43|u0|auto_generated|dffe2~q ),
	.dffe31(\u43|u0|auto_generated|dffe3~q ),
	.dffe41(\u43|u0|auto_generated|dffe4~q ),
	.dffe51(\u43|u0|auto_generated|dffe5~q ),
	.dffe61(\u43|u0|auto_generated|dffe6~q ),
	.dffe71(\u43|u0|auto_generated|dffe7~q ),
	.dffe81(\u43|u0|auto_generated|dffe8~q ),
	.dffe91(\u43|u0|auto_generated|dffe9~q ),
	.dffe101(\u43|u0|auto_generated|dffe10~q ),
	.dffe111(\u43|u0|auto_generated|dffe11~q ),
	.dffe121(\u43|u0|auto_generated|dffe12~q ),
	.dffe131(\u43|u0|auto_generated|dffe13~q ),
	.dffe141(\u43|u0|auto_generated|dffe14~q ),
	.dffe151(\u43|u0|auto_generated|dffe15~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_cordic_sxor_1p_lpm_14 u49(
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.dffe18(\u49|u0|auto_generated|dffe18~q ),
	.dffe1(\u49|u0|auto_generated|dffe1~q ),
	.dffe2(\u49|u0|auto_generated|dffe2~q ),
	.dffe3(\u49|u0|auto_generated|dffe3~q ),
	.dffe4(\u49|u0|auto_generated|dffe4~q ),
	.dffe5(\u49|u0|auto_generated|dffe5~q ),
	.dffe6(\u49|u0|auto_generated|dffe6~q ),
	.dffe7(\u49|u0|auto_generated|dffe7~q ),
	.dffe8(\u49|u0|auto_generated|dffe8~q ),
	.dffe9(\u49|u0|auto_generated|dffe9~q ),
	.dffe10(\u49|u0|auto_generated|dffe10~q ),
	.dffe11(\u49|u0|auto_generated|dffe11~q ),
	.dffe12(\u49|u0|auto_generated|dffe12~q ),
	.dffe13(\u49|u0|auto_generated|dffe13~q ),
	.dffe14(\u49|u0|auto_generated|dffe14~q ),
	.dffe15(\u49|u0|auto_generated|dffe15~q ),
	.dffe16(\u49|u0|auto_generated|dffe16~q ),
	.dffe17(\u49|u0|auto_generated|dffe17~q ),
	.dffe161(\u48|u0|auto_generated|dffe16~q ),
	.pipeline_dffe_17(\u47|u0|auto_generated|pipeline_dffe[17]~q ),
	.dffe181(\u46|u0|auto_generated|dffe18~q ),
	.dffe171(\u46|u0|auto_generated|dffe17~q ),
	.pipeline_dffe_16(\u47|u0|auto_generated|pipeline_dffe[16]~q ),
	.dffe19(\u46|u0|auto_generated|dffe1~q ),
	.dffe21(\u46|u0|auto_generated|dffe2~q ),
	.dffe31(\u46|u0|auto_generated|dffe3~q ),
	.dffe41(\u46|u0|auto_generated|dffe4~q ),
	.dffe51(\u46|u0|auto_generated|dffe5~q ),
	.dffe61(\u46|u0|auto_generated|dffe6~q ),
	.dffe71(\u46|u0|auto_generated|dffe7~q ),
	.dffe81(\u46|u0|auto_generated|dffe8~q ),
	.dffe91(\u46|u0|auto_generated|dffe9~q ),
	.dffe101(\u46|u0|auto_generated|dffe10~q ),
	.dffe111(\u46|u0|auto_generated|dffe11~q ),
	.dffe121(\u46|u0|auto_generated|dffe12~q ),
	.dffe131(\u46|u0|auto_generated|dffe13~q ),
	.dffe141(\u46|u0|auto_generated|dffe14~q ),
	.dffe151(\u46|u0|auto_generated|dffe15~q ),
	.dffe162(\u46|u0|auto_generated|dffe16~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_cordic_zxor_1p_lpm_13 u48(
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.dffe16(\u48|u0|auto_generated|dffe16~q ),
	.dffe15(\u48|u0|auto_generated|dffe15~q ),
	.dffe14(\u48|u0|auto_generated|dffe14~q ),
	.dffe161(\u45|u0|auto_generated|dffe16~q ),
	.dffe13(\u48|u0|auto_generated|dffe13~q ),
	.dffe12(\u48|u0|auto_generated|dffe12~q ),
	.dffe151(\u45|u0|auto_generated|dffe15~q ),
	.dffe11(\u48|u0|auto_generated|dffe11~q ),
	.dffe141(\u45|u0|auto_generated|dffe14~q ),
	.dffe10(\u48|u0|auto_generated|dffe10~q ),
	.dffe131(\u45|u0|auto_generated|dffe13~q ),
	.dffe9(\u48|u0|auto_generated|dffe9~q ),
	.dffe121(\u45|u0|auto_generated|dffe12~q ),
	.dffe8(\u48|u0|auto_generated|dffe8~q ),
	.dffe111(\u45|u0|auto_generated|dffe11~q ),
	.dffe7(\u48|u0|auto_generated|dffe7~q ),
	.dffe101(\u45|u0|auto_generated|dffe10~q ),
	.dffe6(\u48|u0|auto_generated|dffe6~q ),
	.dffe91(\u45|u0|auto_generated|dffe9~q ),
	.dffe5(\u48|u0|auto_generated|dffe5~q ),
	.dffe81(\u45|u0|auto_generated|dffe8~q ),
	.dffe4(\u48|u0|auto_generated|dffe4~q ),
	.dffe71(\u45|u0|auto_generated|dffe7~q ),
	.dffe3(\u48|u0|auto_generated|dffe3~q ),
	.dffe61(\u45|u0|auto_generated|dffe6~q ),
	.dffe2(\u48|u0|auto_generated|dffe2~q ),
	.dffe51(\u45|u0|auto_generated|dffe5~q ),
	.dffe1(\u48|u0|auto_generated|dffe1~q ),
	.dffe41(\u45|u0|auto_generated|dffe4~q ),
	.dffe31(\u45|u0|auto_generated|dffe3~q ),
	.dffe21(\u45|u0|auto_generated|dffe2~q ),
	.dffe17(\u45|u0|auto_generated|dffe1~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_cordic_zxor_1p_lpm_14 u51(
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.dffe16(\u51|u0|auto_generated|dffe16~q ),
	.dffe161(\u48|u0|auto_generated|dffe16~q ),
	.dffe15(\u48|u0|auto_generated|dffe15~q ),
	.dffe14(\u48|u0|auto_generated|dffe14~q ),
	.dffe13(\u48|u0|auto_generated|dffe13~q ),
	.dffe12(\u48|u0|auto_generated|dffe12~q ),
	.dffe11(\u48|u0|auto_generated|dffe11~q ),
	.dffe10(\u48|u0|auto_generated|dffe10~q ),
	.dffe9(\u48|u0|auto_generated|dffe9~q ),
	.dffe8(\u48|u0|auto_generated|dffe8~q ),
	.dffe7(\u48|u0|auto_generated|dffe7~q ),
	.dffe6(\u48|u0|auto_generated|dffe6~q ),
	.dffe5(\u48|u0|auto_generated|dffe5~q ),
	.dffe4(\u48|u0|auto_generated|dffe4~q ),
	.dffe3(\u48|u0|auto_generated|dffe3~q ),
	.dffe2(\u48|u0|auto_generated|dffe2~q ),
	.dffe1(\u48|u0|auto_generated|dffe1~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_cordic_axor_1p_lpm_14 u50(
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.pipeline_dffe_17(\u50|u0|auto_generated|pipeline_dffe[17]~q ),
	.pipeline_dffe_0(\u50|u0|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_1(\u50|u0|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_2(\u50|u0|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\u50|u0|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\u50|u0|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\u50|u0|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\u50|u0|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\u50|u0|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\u50|u0|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\u50|u0|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_10(\u50|u0|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_11(\u50|u0|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_12(\u50|u0|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_13(\u50|u0|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_14(\u50|u0|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_15(\u50|u0|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_16(\u50|u0|auto_generated|pipeline_dffe[16]~q ),
	.dffe16(\u48|u0|auto_generated|dffe16~q ),
	.pipeline_dffe_171(\u47|u0|auto_generated|pipeline_dffe[17]~q ),
	.dffe18(\u46|u0|auto_generated|dffe18~q ),
	.dffe17(\u46|u0|auto_generated|dffe17~q ),
	.pipeline_dffe_161(\u47|u0|auto_generated|pipeline_dffe[16]~q ),
	.pipeline_dffe_01(\u47|u0|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_18(\u47|u0|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_21(\u47|u0|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_31(\u47|u0|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_41(\u47|u0|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_51(\u47|u0|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_61(\u47|u0|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_71(\u47|u0|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_81(\u47|u0|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_91(\u47|u0|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_101(\u47|u0|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_111(\u47|u0|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_121(\u47|u0|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_131(\u47|u0|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_141(\u47|u0|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_151(\u47|u0|auto_generated|pipeline_dffe[15]~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_cordic_axor_1p_lpm_15 u53(
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.pipeline_dffe_0(\u53|u0|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_1(\u53|u0|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_2(\u53|u0|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\u53|u0|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\u53|u0|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\u53|u0|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\u53|u0|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\u53|u0|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\u53|u0|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\u53|u0|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_10(\u53|u0|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_11(\u53|u0|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_12(\u53|u0|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_13(\u53|u0|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_14(\u53|u0|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_15(\u53|u0|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_16(\u53|u0|auto_generated|pipeline_dffe[16]~q ),
	.pipeline_dffe_17(\u53|u0|auto_generated|pipeline_dffe[17]~q ),
	.dffe16(\u51|u0|auto_generated|dffe16~q ),
	.dffe18(\u49|u0|auto_generated|dffe18~q ),
	.pipeline_dffe_171(\u50|u0|auto_generated|pipeline_dffe[17]~q ),
	.pipeline_dffe_01(\u50|u0|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_18(\u50|u0|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_21(\u50|u0|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_31(\u50|u0|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_41(\u50|u0|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_51(\u50|u0|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_61(\u50|u0|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_71(\u50|u0|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_81(\u50|u0|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_91(\u50|u0|auto_generated|pipeline_dffe[9]~q ),
	.pipeline_dffe_101(\u50|u0|auto_generated|pipeline_dffe[10]~q ),
	.pipeline_dffe_111(\u50|u0|auto_generated|pipeline_dffe[11]~q ),
	.pipeline_dffe_121(\u50|u0|auto_generated|pipeline_dffe[12]~q ),
	.pipeline_dffe_131(\u50|u0|auto_generated|pipeline_dffe[13]~q ),
	.pipeline_dffe_141(\u50|u0|auto_generated|pipeline_dffe[14]~q ),
	.pipeline_dffe_151(\u50|u0|auto_generated|pipeline_dffe[15]~q ),
	.pipeline_dffe_161(\u50|u0|auto_generated|pipeline_dffe[16]~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_cordic_sxor_1p_lpm_15 u52(
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.dffe1(\u52|u0|auto_generated|dffe1~q ),
	.dffe2(\u52|u0|auto_generated|dffe2~q ),
	.dffe3(\u52|u0|auto_generated|dffe3~q ),
	.dffe4(\u52|u0|auto_generated|dffe4~q ),
	.dffe5(\u52|u0|auto_generated|dffe5~q ),
	.dffe6(\u52|u0|auto_generated|dffe6~q ),
	.dffe7(\u52|u0|auto_generated|dffe7~q ),
	.dffe8(\u52|u0|auto_generated|dffe8~q ),
	.dffe9(\u52|u0|auto_generated|dffe9~q ),
	.dffe10(\u52|u0|auto_generated|dffe10~q ),
	.dffe11(\u52|u0|auto_generated|dffe11~q ),
	.dffe12(\u52|u0|auto_generated|dffe12~q ),
	.dffe13(\u52|u0|auto_generated|dffe13~q ),
	.dffe14(\u52|u0|auto_generated|dffe14~q ),
	.dffe15(\u52|u0|auto_generated|dffe15~q ),
	.dffe16(\u52|u0|auto_generated|dffe16~q ),
	.dffe17(\u52|u0|auto_generated|dffe17~q ),
	.dffe18(\u52|u0|auto_generated|dffe18~q ),
	.dffe161(\u51|u0|auto_generated|dffe16~q ),
	.dffe181(\u49|u0|auto_generated|dffe18~q ),
	.pipeline_dffe_17(\u50|u0|auto_generated|pipeline_dffe[17]~q ),
	.dffe19(\u49|u0|auto_generated|dffe1~q ),
	.dffe21(\u49|u0|auto_generated|dffe2~q ),
	.dffe31(\u49|u0|auto_generated|dffe3~q ),
	.dffe41(\u49|u0|auto_generated|dffe4~q ),
	.dffe51(\u49|u0|auto_generated|dffe5~q ),
	.dffe61(\u49|u0|auto_generated|dffe6~q ),
	.dffe71(\u49|u0|auto_generated|dffe7~q ),
	.dffe81(\u49|u0|auto_generated|dffe8~q ),
	.dffe91(\u49|u0|auto_generated|dffe9~q ),
	.dffe101(\u49|u0|auto_generated|dffe10~q ),
	.dffe111(\u49|u0|auto_generated|dffe11~q ),
	.dffe121(\u49|u0|auto_generated|dffe12~q ),
	.dffe131(\u49|u0|auto_generated|dffe13~q ),
	.dffe141(\u49|u0|auto_generated|dffe14~q ),
	.dffe151(\u49|u0|auto_generated|dffe15~q ),
	.dffe162(\u49|u0|auto_generated|dffe16~q ),
	.dffe171(\u49|u0|auto_generated|dffe17~q ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_asj_nco_isdr ux710isdr(
	.data_ready1(data_ready),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_dop_reg dop(
	.sin_o_0(sin_o_0),
	.sin_o_1(sin_o_1),
	.sin_o_2(sin_o_2),
	.sin_o_3(sin_o_3),
	.sin_o_4(sin_o_4),
	.sin_o_5(sin_o_5),
	.sin_o_6(sin_o_6),
	.sin_o_7(sin_o_7),
	.sin_o_8(sin_o_8),
	.sin_o_9(sin_o_9),
	.sin_o_10(sin_o_10),
	.sin_o_11(sin_o_11),
	.sin_o_12(sin_o_12),
	.sin_o_13(sin_o_13),
	.sin_o_14(sin_o_14),
	.sin_o_15(sin_o_15),
	.sin_o_16(sin_o_16),
	.sin_o_17(sin_o_17),
	.cos_o_0(cos_o_0),
	.cos_o_1(cos_o_1),
	.cos_o_2(cos_o_2),
	.cos_o_3(cos_o_3),
	.cos_o_4(cos_o_4),
	.cos_o_5(cos_o_5),
	.cos_o_6(cos_o_6),
	.cos_o_7(cos_o_7),
	.cos_o_8(cos_o_8),
	.cos_o_9(cos_o_9),
	.cos_o_10(cos_o_10),
	.cos_o_11(cos_o_11),
	.cos_o_12(cos_o_12),
	.cos_o_13(cos_o_13),
	.cos_o_14(cos_o_14),
	.cos_o_15(cos_o_15),
	.cos_o_16(cos_o_16),
	.cos_o_17(cos_o_17),
	.sin_o_01(\ux005|sin_o[0]~q ),
	.sin_o_18(\ux005|sin_o[1]~q ),
	.sin_o_21(\ux005|sin_o[2]~q ),
	.sin_o_31(\ux005|sin_o[3]~q ),
	.sin_o_41(\ux005|sin_o[4]~q ),
	.sin_o_51(\ux005|sin_o[5]~q ),
	.sin_o_61(\ux005|sin_o[6]~q ),
	.sin_o_71(\ux005|sin_o[7]~q ),
	.sin_o_81(\ux005|sin_o[8]~q ),
	.sin_o_91(\ux005|sin_o[9]~q ),
	.sin_o_101(\ux005|sin_o[10]~q ),
	.sin_o_111(\ux005|sin_o[11]~q ),
	.sin_o_121(\ux005|sin_o[12]~q ),
	.sin_o_131(\ux005|sin_o[13]~q ),
	.sin_o_141(\ux005|sin_o[14]~q ),
	.sin_o_151(\ux005|sin_o[15]~q ),
	.sin_o_161(\ux005|sin_o[16]~q ),
	.sin_o_171(\ux005|sin_o[17]~q ),
	.cos_o_01(\ux005|cos_o[0]~q ),
	.cos_o_18(\ux005|cos_o[1]~q ),
	.cos_o_21(\ux005|cos_o[2]~q ),
	.cos_o_31(\ux005|cos_o[3]~q ),
	.cos_o_41(\ux005|cos_o[4]~q ),
	.cos_o_51(\ux005|cos_o[5]~q ),
	.cos_o_61(\ux005|cos_o[6]~q ),
	.cos_o_71(\ux005|cos_o[7]~q ),
	.cos_o_81(\ux005|cos_o[8]~q ),
	.cos_o_91(\ux005|cos_o[9]~q ),
	.cos_o_101(\ux005|cos_o[10]~q ),
	.cos_o_111(\ux005|cos_o[11]~q ),
	.cos_o_121(\ux005|cos_o[12]~q ),
	.cos_o_131(\ux005|cos_o[13]~q ),
	.cos_o_141(\ux005|cos_o[14]~q ),
	.cos_o_151(\ux005|cos_o[15]~q ),
	.cos_o_161(\ux005|cos_o[16]~q ),
	.cos_o_171(\ux005|cos_o[17]~q ),
	.sin_o_02(\dop|sin_o[0]~0_combout ),
	.clk(clk),
	.reset_n(reset_n),
	.clken(clken));

nco_test_asj_crd_par ux005(
	.sin_o_0(\ux005|sin_o[0]~q ),
	.sin_o_1(\ux005|sin_o[1]~q ),
	.sin_o_2(\ux005|sin_o[2]~q ),
	.sin_o_3(\ux005|sin_o[3]~q ),
	.sin_o_4(\ux005|sin_o[4]~q ),
	.sin_o_5(\ux005|sin_o[5]~q ),
	.sin_o_6(\ux005|sin_o[6]~q ),
	.sin_o_7(\ux005|sin_o[7]~q ),
	.sin_o_8(\ux005|sin_o[8]~q ),
	.sin_o_9(\ux005|sin_o[9]~q ),
	.sin_o_10(\ux005|sin_o[10]~q ),
	.sin_o_11(\ux005|sin_o[11]~q ),
	.sin_o_12(\ux005|sin_o[12]~q ),
	.sin_o_13(\ux005|sin_o[13]~q ),
	.sin_o_14(\ux005|sin_o[14]~q ),
	.sin_o_15(\ux005|sin_o[15]~q ),
	.sin_o_16(\ux005|sin_o[16]~q ),
	.sin_o_17(\ux005|sin_o[17]~q ),
	.cos_o_0(\ux005|cos_o[0]~q ),
	.cos_o_1(\ux005|cos_o[1]~q ),
	.cos_o_2(\ux005|cos_o[2]~q ),
	.cos_o_3(\ux005|cos_o[3]~q ),
	.cos_o_4(\ux005|cos_o[4]~q ),
	.cos_o_5(\ux005|cos_o[5]~q ),
	.cos_o_6(\ux005|cos_o[6]~q ),
	.cos_o_7(\ux005|cos_o[7]~q ),
	.cos_o_8(\ux005|cos_o[8]~q ),
	.cos_o_9(\ux005|cos_o[9]~q ),
	.cos_o_10(\ux005|cos_o[10]~q ),
	.cos_o_11(\ux005|cos_o[11]~q ),
	.cos_o_12(\ux005|cos_o[12]~q ),
	.cos_o_13(\ux005|cos_o[13]~q ),
	.cos_o_14(\ux005|cos_o[14]~q ),
	.cos_o_15(\ux005|cos_o[15]~q ),
	.cos_o_16(\ux005|cos_o[16]~q ),
	.cos_o_17(\ux005|cos_o[17]~q ),
	.cordic_y_res_d_0(\cordinv|cordic_y_res_d[0]~q ),
	.cordic_y_res_2c_0(\cordinv|cordic_y_res_2c[0]~q ),
	.cordic_x_res_d_0(\cordinv|cordic_x_res_d[0]~q ),
	.cordic_x_res_2c_0(\cordinv|cordic_x_res_2c[0]~q ),
	.seg_rot_1(\css|seg_rot[1]~q ),
	.seg_rot_0(\css|seg_rot[0]~q ),
	.cordic_y_res_d_1(\cordinv|cordic_y_res_d[1]~q ),
	.cordic_y_res_2c_1(\cordinv|cordic_y_res_2c[1]~q ),
	.cordic_x_res_d_1(\cordinv|cordic_x_res_d[1]~q ),
	.cordic_x_res_2c_1(\cordinv|cordic_x_res_2c[1]~q ),
	.cordic_y_res_d_2(\cordinv|cordic_y_res_d[2]~q ),
	.cordic_y_res_2c_2(\cordinv|cordic_y_res_2c[2]~q ),
	.cordic_x_res_d_2(\cordinv|cordic_x_res_d[2]~q ),
	.cordic_x_res_2c_2(\cordinv|cordic_x_res_2c[2]~q ),
	.cordic_y_res_d_3(\cordinv|cordic_y_res_d[3]~q ),
	.cordic_y_res_2c_3(\cordinv|cordic_y_res_2c[3]~q ),
	.cordic_x_res_d_3(\cordinv|cordic_x_res_d[3]~q ),
	.cordic_x_res_2c_3(\cordinv|cordic_x_res_2c[3]~q ),
	.cordic_y_res_d_4(\cordinv|cordic_y_res_d[4]~q ),
	.cordic_y_res_2c_4(\cordinv|cordic_y_res_2c[4]~q ),
	.cordic_x_res_d_4(\cordinv|cordic_x_res_d[4]~q ),
	.cordic_x_res_2c_4(\cordinv|cordic_x_res_2c[4]~q ),
	.cordic_y_res_d_5(\cordinv|cordic_y_res_d[5]~q ),
	.cordic_y_res_2c_5(\cordinv|cordic_y_res_2c[5]~q ),
	.cordic_x_res_d_5(\cordinv|cordic_x_res_d[5]~q ),
	.cordic_x_res_2c_5(\cordinv|cordic_x_res_2c[5]~q ),
	.cordic_y_res_d_6(\cordinv|cordic_y_res_d[6]~q ),
	.cordic_y_res_2c_6(\cordinv|cordic_y_res_2c[6]~q ),
	.cordic_x_res_d_6(\cordinv|cordic_x_res_d[6]~q ),
	.cordic_x_res_2c_6(\cordinv|cordic_x_res_2c[6]~q ),
	.cordic_y_res_d_7(\cordinv|cordic_y_res_d[7]~q ),
	.cordic_y_res_2c_7(\cordinv|cordic_y_res_2c[7]~q ),
	.cordic_x_res_d_7(\cordinv|cordic_x_res_d[7]~q ),
	.cordic_x_res_2c_7(\cordinv|cordic_x_res_2c[7]~q ),
	.cordic_y_res_d_8(\cordinv|cordic_y_res_d[8]~q ),
	.cordic_y_res_2c_8(\cordinv|cordic_y_res_2c[8]~q ),
	.cordic_x_res_d_8(\cordinv|cordic_x_res_d[8]~q ),
	.cordic_x_res_2c_8(\cordinv|cordic_x_res_2c[8]~q ),
	.cordic_y_res_d_9(\cordinv|cordic_y_res_d[9]~q ),
	.cordic_y_res_2c_9(\cordinv|cordic_y_res_2c[9]~q ),
	.cordic_x_res_d_9(\cordinv|cordic_x_res_d[9]~q ),
	.cordic_x_res_2c_9(\cordinv|cordic_x_res_2c[9]~q ),
	.cordic_y_res_d_10(\cordinv|cordic_y_res_d[10]~q ),
	.cordic_y_res_2c_10(\cordinv|cordic_y_res_2c[10]~q ),
	.cordic_x_res_d_10(\cordinv|cordic_x_res_d[10]~q ),
	.cordic_x_res_2c_10(\cordinv|cordic_x_res_2c[10]~q ),
	.cordic_y_res_d_11(\cordinv|cordic_y_res_d[11]~q ),
	.cordic_y_res_2c_11(\cordinv|cordic_y_res_2c[11]~q ),
	.cordic_x_res_d_11(\cordinv|cordic_x_res_d[11]~q ),
	.cordic_x_res_2c_11(\cordinv|cordic_x_res_2c[11]~q ),
	.cordic_y_res_d_12(\cordinv|cordic_y_res_d[12]~q ),
	.cordic_y_res_2c_12(\cordinv|cordic_y_res_2c[12]~q ),
	.cordic_x_res_d_12(\cordinv|cordic_x_res_d[12]~q ),
	.cordic_x_res_2c_12(\cordinv|cordic_x_res_2c[12]~q ),
	.cordic_y_res_d_13(\cordinv|cordic_y_res_d[13]~q ),
	.cordic_y_res_2c_13(\cordinv|cordic_y_res_2c[13]~q ),
	.cordic_x_res_d_13(\cordinv|cordic_x_res_d[13]~q ),
	.cordic_x_res_2c_13(\cordinv|cordic_x_res_2c[13]~q ),
	.cordic_y_res_d_14(\cordinv|cordic_y_res_d[14]~q ),
	.cordic_y_res_2c_14(\cordinv|cordic_y_res_2c[14]~q ),
	.cordic_x_res_d_14(\cordinv|cordic_x_res_d[14]~q ),
	.cordic_x_res_2c_14(\cordinv|cordic_x_res_2c[14]~q ),
	.cordic_y_res_d_15(\cordinv|cordic_y_res_d[15]~q ),
	.cordic_y_res_2c_15(\cordinv|cordic_y_res_2c[15]~q ),
	.cordic_x_res_d_15(\cordinv|cordic_x_res_d[15]~q ),
	.cordic_x_res_2c_15(\cordinv|cordic_x_res_2c[15]~q ),
	.cordic_y_res_d_16(\cordinv|cordic_y_res_d[16]~q ),
	.cordic_y_res_2c_16(\cordinv|cordic_y_res_2c[16]~q ),
	.cordic_x_res_d_16(\cordinv|cordic_x_res_d[16]~q ),
	.cordic_x_res_2c_16(\cordinv|cordic_x_res_2c[16]~q ),
	.cordic_y_res_d_17(\cordinv|cordic_y_res_d[17]~q ),
	.cordic_y_res_2c_17(\cordinv|cordic_y_res_2c[17]~q ),
	.cordic_x_res_d_17(\cordinv|cordic_x_res_d[17]~q ),
	.cordic_x_res_2c_17(\cordinv|cordic_x_res_2c[17]~q ),
	.sin_o_01(\dop|sin_o[0]~0_combout ),
	.clk(clk),
	.reset_n(reset_n));

nco_test_cord_2c cordinv(
	.cordic_y_res_d_0(\cordinv|cordic_y_res_d[0]~q ),
	.cordic_y_res_2c_0(\cordinv|cordic_y_res_2c[0]~q ),
	.cordic_x_res_d_0(\cordinv|cordic_x_res_d[0]~q ),
	.cordic_x_res_2c_0(\cordinv|cordic_x_res_2c[0]~q ),
	.cordic_y_res_d_1(\cordinv|cordic_y_res_d[1]~q ),
	.cordic_y_res_2c_1(\cordinv|cordic_y_res_2c[1]~q ),
	.cordic_x_res_d_1(\cordinv|cordic_x_res_d[1]~q ),
	.cordic_x_res_2c_1(\cordinv|cordic_x_res_2c[1]~q ),
	.cordic_y_res_d_2(\cordinv|cordic_y_res_d[2]~q ),
	.cordic_y_res_2c_2(\cordinv|cordic_y_res_2c[2]~q ),
	.cordic_x_res_d_2(\cordinv|cordic_x_res_d[2]~q ),
	.cordic_x_res_2c_2(\cordinv|cordic_x_res_2c[2]~q ),
	.cordic_y_res_d_3(\cordinv|cordic_y_res_d[3]~q ),
	.cordic_y_res_2c_3(\cordinv|cordic_y_res_2c[3]~q ),
	.cordic_x_res_d_3(\cordinv|cordic_x_res_d[3]~q ),
	.cordic_x_res_2c_3(\cordinv|cordic_x_res_2c[3]~q ),
	.cordic_y_res_d_4(\cordinv|cordic_y_res_d[4]~q ),
	.cordic_y_res_2c_4(\cordinv|cordic_y_res_2c[4]~q ),
	.cordic_x_res_d_4(\cordinv|cordic_x_res_d[4]~q ),
	.cordic_x_res_2c_4(\cordinv|cordic_x_res_2c[4]~q ),
	.cordic_y_res_d_5(\cordinv|cordic_y_res_d[5]~q ),
	.cordic_y_res_2c_5(\cordinv|cordic_y_res_2c[5]~q ),
	.cordic_x_res_d_5(\cordinv|cordic_x_res_d[5]~q ),
	.cordic_x_res_2c_5(\cordinv|cordic_x_res_2c[5]~q ),
	.cordic_y_res_d_6(\cordinv|cordic_y_res_d[6]~q ),
	.cordic_y_res_2c_6(\cordinv|cordic_y_res_2c[6]~q ),
	.cordic_x_res_d_6(\cordinv|cordic_x_res_d[6]~q ),
	.cordic_x_res_2c_6(\cordinv|cordic_x_res_2c[6]~q ),
	.cordic_y_res_d_7(\cordinv|cordic_y_res_d[7]~q ),
	.cordic_y_res_2c_7(\cordinv|cordic_y_res_2c[7]~q ),
	.cordic_x_res_d_7(\cordinv|cordic_x_res_d[7]~q ),
	.cordic_x_res_2c_7(\cordinv|cordic_x_res_2c[7]~q ),
	.cordic_y_res_d_8(\cordinv|cordic_y_res_d[8]~q ),
	.cordic_y_res_2c_8(\cordinv|cordic_y_res_2c[8]~q ),
	.cordic_x_res_d_8(\cordinv|cordic_x_res_d[8]~q ),
	.cordic_x_res_2c_8(\cordinv|cordic_x_res_2c[8]~q ),
	.cordic_y_res_d_9(\cordinv|cordic_y_res_d[9]~q ),
	.cordic_y_res_2c_9(\cordinv|cordic_y_res_2c[9]~q ),
	.cordic_x_res_d_9(\cordinv|cordic_x_res_d[9]~q ),
	.cordic_x_res_2c_9(\cordinv|cordic_x_res_2c[9]~q ),
	.cordic_y_res_d_10(\cordinv|cordic_y_res_d[10]~q ),
	.cordic_y_res_2c_10(\cordinv|cordic_y_res_2c[10]~q ),
	.cordic_x_res_d_10(\cordinv|cordic_x_res_d[10]~q ),
	.cordic_x_res_2c_10(\cordinv|cordic_x_res_2c[10]~q ),
	.cordic_y_res_d_11(\cordinv|cordic_y_res_d[11]~q ),
	.cordic_y_res_2c_11(\cordinv|cordic_y_res_2c[11]~q ),
	.cordic_x_res_d_11(\cordinv|cordic_x_res_d[11]~q ),
	.cordic_x_res_2c_11(\cordinv|cordic_x_res_2c[11]~q ),
	.cordic_y_res_d_12(\cordinv|cordic_y_res_d[12]~q ),
	.cordic_y_res_2c_12(\cordinv|cordic_y_res_2c[12]~q ),
	.cordic_x_res_d_12(\cordinv|cordic_x_res_d[12]~q ),
	.cordic_x_res_2c_12(\cordinv|cordic_x_res_2c[12]~q ),
	.cordic_y_res_d_13(\cordinv|cordic_y_res_d[13]~q ),
	.cordic_y_res_2c_13(\cordinv|cordic_y_res_2c[13]~q ),
	.cordic_x_res_d_13(\cordinv|cordic_x_res_d[13]~q ),
	.cordic_x_res_2c_13(\cordinv|cordic_x_res_2c[13]~q ),
	.cordic_y_res_d_14(\cordinv|cordic_y_res_d[14]~q ),
	.cordic_y_res_2c_14(\cordinv|cordic_y_res_2c[14]~q ),
	.cordic_x_res_d_14(\cordinv|cordic_x_res_d[14]~q ),
	.cordic_x_res_2c_14(\cordinv|cordic_x_res_2c[14]~q ),
	.cordic_y_res_d_15(\cordinv|cordic_y_res_d[15]~q ),
	.cordic_y_res_2c_15(\cordinv|cordic_y_res_2c[15]~q ),
	.cordic_x_res_d_15(\cordinv|cordic_x_res_d[15]~q ),
	.cordic_x_res_2c_15(\cordinv|cordic_x_res_2c[15]~q ),
	.cordic_y_res_d_16(\cordinv|cordic_y_res_d[16]~q ),
	.cordic_y_res_2c_16(\cordinv|cordic_y_res_2c[16]~q ),
	.cordic_x_res_d_16(\cordinv|cordic_x_res_d[16]~q ),
	.cordic_x_res_2c_16(\cordinv|cordic_x_res_2c[16]~q ),
	.cordic_y_res_d_17(\cordinv|cordic_y_res_d[17]~q ),
	.cordic_y_res_2c_17(\cordinv|cordic_y_res_2c[17]~q ),
	.cordic_x_res_d_17(\cordinv|cordic_x_res_d[17]~q ),
	.cordic_x_res_2c_17(\cordinv|cordic_x_res_2c[17]~q ),
	.sin_o_0(\dop|sin_o[0]~0_combout ),
	.pipeline_dffe_0(\u53|u0|auto_generated|pipeline_dffe[0]~q ),
	.dffe1(\u52|u0|auto_generated|dffe1~q ),
	.pipeline_dffe_1(\u53|u0|auto_generated|pipeline_dffe[1]~q ),
	.dffe2(\u52|u0|auto_generated|dffe2~q ),
	.pipeline_dffe_2(\u53|u0|auto_generated|pipeline_dffe[2]~q ),
	.dffe3(\u52|u0|auto_generated|dffe3~q ),
	.pipeline_dffe_3(\u53|u0|auto_generated|pipeline_dffe[3]~q ),
	.dffe4(\u52|u0|auto_generated|dffe4~q ),
	.pipeline_dffe_4(\u53|u0|auto_generated|pipeline_dffe[4]~q ),
	.dffe5(\u52|u0|auto_generated|dffe5~q ),
	.pipeline_dffe_5(\u53|u0|auto_generated|pipeline_dffe[5]~q ),
	.dffe6(\u52|u0|auto_generated|dffe6~q ),
	.pipeline_dffe_6(\u53|u0|auto_generated|pipeline_dffe[6]~q ),
	.dffe7(\u52|u0|auto_generated|dffe7~q ),
	.pipeline_dffe_7(\u53|u0|auto_generated|pipeline_dffe[7]~q ),
	.dffe8(\u52|u0|auto_generated|dffe8~q ),
	.pipeline_dffe_8(\u53|u0|auto_generated|pipeline_dffe[8]~q ),
	.dffe9(\u52|u0|auto_generated|dffe9~q ),
	.pipeline_dffe_9(\u53|u0|auto_generated|pipeline_dffe[9]~q ),
	.dffe10(\u52|u0|auto_generated|dffe10~q ),
	.pipeline_dffe_10(\u53|u0|auto_generated|pipeline_dffe[10]~q ),
	.dffe11(\u52|u0|auto_generated|dffe11~q ),
	.pipeline_dffe_11(\u53|u0|auto_generated|pipeline_dffe[11]~q ),
	.dffe12(\u52|u0|auto_generated|dffe12~q ),
	.pipeline_dffe_12(\u53|u0|auto_generated|pipeline_dffe[12]~q ),
	.dffe13(\u52|u0|auto_generated|dffe13~q ),
	.pipeline_dffe_13(\u53|u0|auto_generated|pipeline_dffe[13]~q ),
	.dffe14(\u52|u0|auto_generated|dffe14~q ),
	.pipeline_dffe_14(\u53|u0|auto_generated|pipeline_dffe[14]~q ),
	.dffe15(\u52|u0|auto_generated|dffe15~q ),
	.pipeline_dffe_15(\u53|u0|auto_generated|pipeline_dffe[15]~q ),
	.dffe16(\u52|u0|auto_generated|dffe16~q ),
	.pipeline_dffe_16(\u53|u0|auto_generated|pipeline_dffe[16]~q ),
	.dffe17(\u52|u0|auto_generated|dffe17~q ),
	.pipeline_dffe_17(\u53|u0|auto_generated|pipeline_dffe[17]~q ),
	.dffe18(\u52|u0|auto_generated|dffe18~q ),
	.clk(clk),
	.reset_n(reset_n));

endmodule

module nco_test_asj_altqmcpipe (
	sin_o_0,
	pipeline_dffe_31,
	pipeline_dffe_30,
	pipeline_dffe_29,
	pipeline_dffe_28,
	pipeline_dffe_27,
	pipeline_dffe_26,
	pipeline_dffe_25,
	pipeline_dffe_24,
	pipeline_dffe_23,
	pipeline_dffe_22,
	pipeline_dffe_21,
	pipeline_dffe_20,
	pipeline_dffe_19,
	pipeline_dffe_18,
	pipeline_dffe_17,
	pipeline_dffe_16,
	pipeline_dffe_15,
	pipeline_dffe_14,
	pipeline_dffe_13,
	pipeline_dffe_12,
	pipeline_dffe_11,
	clk,
	reset_n,
	clken,
	phi_inc_i_31,
	phi_inc_i_30,
	phi_inc_i_29,
	phi_inc_i_28,
	phi_inc_i_27,
	phi_inc_i_26,
	phi_inc_i_25,
	phi_inc_i_24,
	phi_inc_i_23,
	phi_inc_i_22,
	phi_inc_i_21,
	phi_inc_i_20,
	phi_inc_i_19,
	phi_inc_i_18,
	phi_inc_i_17,
	phi_inc_i_16,
	phi_inc_i_15,
	phi_inc_i_14,
	phi_inc_i_13,
	phi_inc_i_12,
	phi_inc_i_11,
	phi_inc_i_10,
	phi_inc_i_9,
	phi_inc_i_8,
	phi_inc_i_7,
	phi_inc_i_6,
	phi_inc_i_5,
	phi_inc_i_4,
	phi_inc_i_3,
	phi_inc_i_2,
	phi_inc_i_1,
	phi_inc_i_0)/* synthesis synthesis_greybox=1 */;
input 	sin_o_0;
output 	pipeline_dffe_31;
output 	pipeline_dffe_30;
output 	pipeline_dffe_29;
output 	pipeline_dffe_28;
output 	pipeline_dffe_27;
output 	pipeline_dffe_26;
output 	pipeline_dffe_25;
output 	pipeline_dffe_24;
output 	pipeline_dffe_23;
output 	pipeline_dffe_22;
output 	pipeline_dffe_21;
output 	pipeline_dffe_20;
output 	pipeline_dffe_19;
output 	pipeline_dffe_18;
output 	pipeline_dffe_17;
output 	pipeline_dffe_16;
output 	pipeline_dffe_15;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
input 	clk;
input 	reset_n;
input 	clken;
input 	phi_inc_i_31;
input 	phi_inc_i_30;
input 	phi_inc_i_29;
input 	phi_inc_i_28;
input 	phi_inc_i_27;
input 	phi_inc_i_26;
input 	phi_inc_i_25;
input 	phi_inc_i_24;
input 	phi_inc_i_23;
input 	phi_inc_i_22;
input 	phi_inc_i_21;
input 	phi_inc_i_20;
input 	phi_inc_i_19;
input 	phi_inc_i_18;
input 	phi_inc_i_17;
input 	phi_inc_i_16;
input 	phi_inc_i_15;
input 	phi_inc_i_14;
input 	phi_inc_i_13;
input 	phi_inc_i_12;
input 	phi_inc_i_11;
input 	phi_inc_i_10;
input 	phi_inc_i_9;
input 	phi_inc_i_8;
input 	phi_inc_i_7;
input 	phi_inc_i_6;
input 	phi_inc_i_5;
input 	phi_inc_i_4;
input 	phi_inc_i_3;
input 	phi_inc_i_2;
input 	phi_inc_i_1;
input 	phi_inc_i_0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \phi_int_arr_reg[31]~q ;
wire \phi_int_arr_reg[30]~q ;
wire \phi_int_arr_reg[29]~q ;
wire \phi_int_arr_reg[28]~q ;
wire \phi_int_arr_reg[27]~q ;
wire \phi_int_arr_reg[26]~q ;
wire \phi_int_arr_reg[25]~q ;
wire \phi_int_arr_reg[24]~q ;
wire \phi_int_arr_reg[23]~q ;
wire \phi_int_arr_reg[22]~q ;
wire \phi_int_arr_reg[21]~q ;
wire \phi_int_arr_reg[20]~q ;
wire \phi_int_arr_reg[19]~q ;
wire \phi_int_arr_reg[18]~q ;
wire \phi_int_arr_reg[17]~q ;
wire \phi_int_arr_reg[16]~q ;
wire \phi_int_arr_reg[15]~q ;
wire \phi_int_arr_reg[14]~q ;
wire \phi_int_arr_reg[13]~q ;
wire \phi_int_arr_reg[12]~q ;
wire \phi_int_arr_reg[11]~q ;
wire \phi_int_arr_reg[10]~q ;
wire \phi_int_arr_reg[9]~q ;
wire \phi_int_arr_reg[8]~q ;
wire \phi_int_arr_reg[7]~q ;
wire \phi_int_arr_reg[6]~q ;
wire \phi_int_arr_reg[5]~q ;
wire \phi_int_arr_reg[4]~q ;
wire \phi_int_arr_reg[3]~q ;
wire \phi_int_arr_reg[2]~q ;
wire \phi_int_arr_reg[1]~q ;
wire \phi_int_arr_reg[0]~q ;


nco_test_lpm_add_sub_1 acc(
	.phi_int_arr_reg_31(\phi_int_arr_reg[31]~q ),
	.phi_int_arr_reg_30(\phi_int_arr_reg[30]~q ),
	.phi_int_arr_reg_29(\phi_int_arr_reg[29]~q ),
	.phi_int_arr_reg_28(\phi_int_arr_reg[28]~q ),
	.phi_int_arr_reg_27(\phi_int_arr_reg[27]~q ),
	.phi_int_arr_reg_26(\phi_int_arr_reg[26]~q ),
	.phi_int_arr_reg_25(\phi_int_arr_reg[25]~q ),
	.phi_int_arr_reg_24(\phi_int_arr_reg[24]~q ),
	.phi_int_arr_reg_23(\phi_int_arr_reg[23]~q ),
	.phi_int_arr_reg_22(\phi_int_arr_reg[22]~q ),
	.phi_int_arr_reg_21(\phi_int_arr_reg[21]~q ),
	.phi_int_arr_reg_20(\phi_int_arr_reg[20]~q ),
	.phi_int_arr_reg_19(\phi_int_arr_reg[19]~q ),
	.phi_int_arr_reg_18(\phi_int_arr_reg[18]~q ),
	.phi_int_arr_reg_17(\phi_int_arr_reg[17]~q ),
	.phi_int_arr_reg_16(\phi_int_arr_reg[16]~q ),
	.phi_int_arr_reg_15(\phi_int_arr_reg[15]~q ),
	.phi_int_arr_reg_14(\phi_int_arr_reg[14]~q ),
	.phi_int_arr_reg_13(\phi_int_arr_reg[13]~q ),
	.phi_int_arr_reg_12(\phi_int_arr_reg[12]~q ),
	.phi_int_arr_reg_11(\phi_int_arr_reg[11]~q ),
	.phi_int_arr_reg_10(\phi_int_arr_reg[10]~q ),
	.phi_int_arr_reg_9(\phi_int_arr_reg[9]~q ),
	.phi_int_arr_reg_8(\phi_int_arr_reg[8]~q ),
	.phi_int_arr_reg_7(\phi_int_arr_reg[7]~q ),
	.phi_int_arr_reg_6(\phi_int_arr_reg[6]~q ),
	.phi_int_arr_reg_5(\phi_int_arr_reg[5]~q ),
	.phi_int_arr_reg_4(\phi_int_arr_reg[4]~q ),
	.phi_int_arr_reg_3(\phi_int_arr_reg[3]~q ),
	.phi_int_arr_reg_2(\phi_int_arr_reg[2]~q ),
	.phi_int_arr_reg_1(\phi_int_arr_reg[1]~q ),
	.phi_int_arr_reg_0(\phi_int_arr_reg[0]~q ),
	.pipeline_dffe_31(pipeline_dffe_31),
	.pipeline_dffe_30(pipeline_dffe_30),
	.pipeline_dffe_29(pipeline_dffe_29),
	.pipeline_dffe_28(pipeline_dffe_28),
	.pipeline_dffe_27(pipeline_dffe_27),
	.pipeline_dffe_26(pipeline_dffe_26),
	.pipeline_dffe_25(pipeline_dffe_25),
	.pipeline_dffe_24(pipeline_dffe_24),
	.pipeline_dffe_23(pipeline_dffe_23),
	.pipeline_dffe_22(pipeline_dffe_22),
	.pipeline_dffe_21(pipeline_dffe_21),
	.pipeline_dffe_20(pipeline_dffe_20),
	.pipeline_dffe_19(pipeline_dffe_19),
	.pipeline_dffe_18(pipeline_dffe_18),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_11(pipeline_dffe_11),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \phi_int_arr_reg[31] (
	.clk(clk),
	.d(phi_inc_i_31),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\phi_int_arr_reg[31]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[31] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[31] .power_up = "low";

dffeas \phi_int_arr_reg[30] (
	.clk(clk),
	.d(phi_inc_i_30),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\phi_int_arr_reg[30]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[30] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[30] .power_up = "low";

dffeas \phi_int_arr_reg[29] (
	.clk(clk),
	.d(phi_inc_i_29),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\phi_int_arr_reg[29]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[29] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[29] .power_up = "low";

dffeas \phi_int_arr_reg[28] (
	.clk(clk),
	.d(phi_inc_i_28),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\phi_int_arr_reg[28]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[28] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[28] .power_up = "low";

dffeas \phi_int_arr_reg[27] (
	.clk(clk),
	.d(phi_inc_i_27),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\phi_int_arr_reg[27]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[27] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[27] .power_up = "low";

dffeas \phi_int_arr_reg[26] (
	.clk(clk),
	.d(phi_inc_i_26),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\phi_int_arr_reg[26]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[26] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[26] .power_up = "low";

dffeas \phi_int_arr_reg[25] (
	.clk(clk),
	.d(phi_inc_i_25),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\phi_int_arr_reg[25]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[25] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[25] .power_up = "low";

dffeas \phi_int_arr_reg[24] (
	.clk(clk),
	.d(phi_inc_i_24),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\phi_int_arr_reg[24]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[24] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[24] .power_up = "low";

dffeas \phi_int_arr_reg[23] (
	.clk(clk),
	.d(phi_inc_i_23),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\phi_int_arr_reg[23]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[23] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[23] .power_up = "low";

dffeas \phi_int_arr_reg[22] (
	.clk(clk),
	.d(phi_inc_i_22),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\phi_int_arr_reg[22]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[22] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[22] .power_up = "low";

dffeas \phi_int_arr_reg[21] (
	.clk(clk),
	.d(phi_inc_i_21),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\phi_int_arr_reg[21]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[21] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[21] .power_up = "low";

dffeas \phi_int_arr_reg[20] (
	.clk(clk),
	.d(phi_inc_i_20),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\phi_int_arr_reg[20]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[20] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[20] .power_up = "low";

dffeas \phi_int_arr_reg[19] (
	.clk(clk),
	.d(phi_inc_i_19),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\phi_int_arr_reg[19]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[19] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[19] .power_up = "low";

dffeas \phi_int_arr_reg[18] (
	.clk(clk),
	.d(phi_inc_i_18),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\phi_int_arr_reg[18]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[18] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[18] .power_up = "low";

dffeas \phi_int_arr_reg[17] (
	.clk(clk),
	.d(phi_inc_i_17),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\phi_int_arr_reg[17]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[17] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[17] .power_up = "low";

dffeas \phi_int_arr_reg[16] (
	.clk(clk),
	.d(phi_inc_i_16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\phi_int_arr_reg[16]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[16] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[16] .power_up = "low";

dffeas \phi_int_arr_reg[15] (
	.clk(clk),
	.d(phi_inc_i_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\phi_int_arr_reg[15]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[15] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[15] .power_up = "low";

dffeas \phi_int_arr_reg[14] (
	.clk(clk),
	.d(phi_inc_i_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\phi_int_arr_reg[14]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[14] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[14] .power_up = "low";

dffeas \phi_int_arr_reg[13] (
	.clk(clk),
	.d(phi_inc_i_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\phi_int_arr_reg[13]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[13] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[13] .power_up = "low";

dffeas \phi_int_arr_reg[12] (
	.clk(clk),
	.d(phi_inc_i_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\phi_int_arr_reg[12]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[12] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[12] .power_up = "low";

dffeas \phi_int_arr_reg[11] (
	.clk(clk),
	.d(phi_inc_i_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\phi_int_arr_reg[11]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[11] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[11] .power_up = "low";

dffeas \phi_int_arr_reg[10] (
	.clk(clk),
	.d(phi_inc_i_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\phi_int_arr_reg[10]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[10] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[10] .power_up = "low";

dffeas \phi_int_arr_reg[9] (
	.clk(clk),
	.d(phi_inc_i_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\phi_int_arr_reg[9]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[9] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[9] .power_up = "low";

dffeas \phi_int_arr_reg[8] (
	.clk(clk),
	.d(phi_inc_i_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\phi_int_arr_reg[8]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[8] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[8] .power_up = "low";

dffeas \phi_int_arr_reg[7] (
	.clk(clk),
	.d(phi_inc_i_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\phi_int_arr_reg[7]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[7] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[7] .power_up = "low";

dffeas \phi_int_arr_reg[6] (
	.clk(clk),
	.d(phi_inc_i_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\phi_int_arr_reg[6]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[6] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[6] .power_up = "low";

dffeas \phi_int_arr_reg[5] (
	.clk(clk),
	.d(phi_inc_i_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\phi_int_arr_reg[5]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[5] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[5] .power_up = "low";

dffeas \phi_int_arr_reg[4] (
	.clk(clk),
	.d(phi_inc_i_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\phi_int_arr_reg[4]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[4] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[4] .power_up = "low";

dffeas \phi_int_arr_reg[3] (
	.clk(clk),
	.d(phi_inc_i_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\phi_int_arr_reg[3]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[3] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[3] .power_up = "low";

dffeas \phi_int_arr_reg[2] (
	.clk(clk),
	.d(phi_inc_i_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\phi_int_arr_reg[2]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[2] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[2] .power_up = "low";

dffeas \phi_int_arr_reg[1] (
	.clk(clk),
	.d(phi_inc_i_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\phi_int_arr_reg[1]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[1] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[1] .power_up = "low";

dffeas \phi_int_arr_reg[0] (
	.clk(clk),
	.d(phi_inc_i_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\phi_int_arr_reg[0]~q ),
	.prn(vcc));
defparam \phi_int_arr_reg[0] .is_wysiwyg = "true";
defparam \phi_int_arr_reg[0] .power_up = "low";

endmodule

module nco_test_lpm_add_sub_1 (
	phi_int_arr_reg_31,
	phi_int_arr_reg_30,
	phi_int_arr_reg_29,
	phi_int_arr_reg_28,
	phi_int_arr_reg_27,
	phi_int_arr_reg_26,
	phi_int_arr_reg_25,
	phi_int_arr_reg_24,
	phi_int_arr_reg_23,
	phi_int_arr_reg_22,
	phi_int_arr_reg_21,
	phi_int_arr_reg_20,
	phi_int_arr_reg_19,
	phi_int_arr_reg_18,
	phi_int_arr_reg_17,
	phi_int_arr_reg_16,
	phi_int_arr_reg_15,
	phi_int_arr_reg_14,
	phi_int_arr_reg_13,
	phi_int_arr_reg_12,
	phi_int_arr_reg_11,
	phi_int_arr_reg_10,
	phi_int_arr_reg_9,
	phi_int_arr_reg_8,
	phi_int_arr_reg_7,
	phi_int_arr_reg_6,
	phi_int_arr_reg_5,
	phi_int_arr_reg_4,
	phi_int_arr_reg_3,
	phi_int_arr_reg_2,
	phi_int_arr_reg_1,
	phi_int_arr_reg_0,
	pipeline_dffe_31,
	pipeline_dffe_30,
	pipeline_dffe_29,
	pipeline_dffe_28,
	pipeline_dffe_27,
	pipeline_dffe_26,
	pipeline_dffe_25,
	pipeline_dffe_24,
	pipeline_dffe_23,
	pipeline_dffe_22,
	pipeline_dffe_21,
	pipeline_dffe_20,
	pipeline_dffe_19,
	pipeline_dffe_18,
	pipeline_dffe_17,
	pipeline_dffe_16,
	pipeline_dffe_15,
	pipeline_dffe_14,
	pipeline_dffe_13,
	pipeline_dffe_12,
	pipeline_dffe_11,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	phi_int_arr_reg_31;
input 	phi_int_arr_reg_30;
input 	phi_int_arr_reg_29;
input 	phi_int_arr_reg_28;
input 	phi_int_arr_reg_27;
input 	phi_int_arr_reg_26;
input 	phi_int_arr_reg_25;
input 	phi_int_arr_reg_24;
input 	phi_int_arr_reg_23;
input 	phi_int_arr_reg_22;
input 	phi_int_arr_reg_21;
input 	phi_int_arr_reg_20;
input 	phi_int_arr_reg_19;
input 	phi_int_arr_reg_18;
input 	phi_int_arr_reg_17;
input 	phi_int_arr_reg_16;
input 	phi_int_arr_reg_15;
input 	phi_int_arr_reg_14;
input 	phi_int_arr_reg_13;
input 	phi_int_arr_reg_12;
input 	phi_int_arr_reg_11;
input 	phi_int_arr_reg_10;
input 	phi_int_arr_reg_9;
input 	phi_int_arr_reg_8;
input 	phi_int_arr_reg_7;
input 	phi_int_arr_reg_6;
input 	phi_int_arr_reg_5;
input 	phi_int_arr_reg_4;
input 	phi_int_arr_reg_3;
input 	phi_int_arr_reg_2;
input 	phi_int_arr_reg_1;
input 	phi_int_arr_reg_0;
output 	pipeline_dffe_31;
output 	pipeline_dffe_30;
output 	pipeline_dffe_29;
output 	pipeline_dffe_28;
output 	pipeline_dffe_27;
output 	pipeline_dffe_26;
output 	pipeline_dffe_25;
output 	pipeline_dffe_24;
output 	pipeline_dffe_23;
output 	pipeline_dffe_22;
output 	pipeline_dffe_21;
output 	pipeline_dffe_20;
output 	pipeline_dffe_19;
output 	pipeline_dffe_18;
output 	pipeline_dffe_17;
output 	pipeline_dffe_16;
output 	pipeline_dffe_15;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_add_sub_jmh auto_generated(
	.phi_int_arr_reg_31(phi_int_arr_reg_31),
	.phi_int_arr_reg_30(phi_int_arr_reg_30),
	.phi_int_arr_reg_29(phi_int_arr_reg_29),
	.phi_int_arr_reg_28(phi_int_arr_reg_28),
	.phi_int_arr_reg_27(phi_int_arr_reg_27),
	.phi_int_arr_reg_26(phi_int_arr_reg_26),
	.phi_int_arr_reg_25(phi_int_arr_reg_25),
	.phi_int_arr_reg_24(phi_int_arr_reg_24),
	.phi_int_arr_reg_23(phi_int_arr_reg_23),
	.phi_int_arr_reg_22(phi_int_arr_reg_22),
	.phi_int_arr_reg_21(phi_int_arr_reg_21),
	.phi_int_arr_reg_20(phi_int_arr_reg_20),
	.phi_int_arr_reg_19(phi_int_arr_reg_19),
	.phi_int_arr_reg_18(phi_int_arr_reg_18),
	.phi_int_arr_reg_17(phi_int_arr_reg_17),
	.phi_int_arr_reg_16(phi_int_arr_reg_16),
	.phi_int_arr_reg_15(phi_int_arr_reg_15),
	.phi_int_arr_reg_14(phi_int_arr_reg_14),
	.phi_int_arr_reg_13(phi_int_arr_reg_13),
	.phi_int_arr_reg_12(phi_int_arr_reg_12),
	.phi_int_arr_reg_11(phi_int_arr_reg_11),
	.phi_int_arr_reg_10(phi_int_arr_reg_10),
	.phi_int_arr_reg_9(phi_int_arr_reg_9),
	.phi_int_arr_reg_8(phi_int_arr_reg_8),
	.phi_int_arr_reg_7(phi_int_arr_reg_7),
	.phi_int_arr_reg_6(phi_int_arr_reg_6),
	.phi_int_arr_reg_5(phi_int_arr_reg_5),
	.phi_int_arr_reg_4(phi_int_arr_reg_4),
	.phi_int_arr_reg_3(phi_int_arr_reg_3),
	.phi_int_arr_reg_2(phi_int_arr_reg_2),
	.phi_int_arr_reg_1(phi_int_arr_reg_1),
	.phi_int_arr_reg_0(phi_int_arr_reg_0),
	.pipeline_dffe_31(pipeline_dffe_31),
	.pipeline_dffe_30(pipeline_dffe_30),
	.pipeline_dffe_29(pipeline_dffe_29),
	.pipeline_dffe_28(pipeline_dffe_28),
	.pipeline_dffe_27(pipeline_dffe_27),
	.pipeline_dffe_26(pipeline_dffe_26),
	.pipeline_dffe_25(pipeline_dffe_25),
	.pipeline_dffe_24(pipeline_dffe_24),
	.pipeline_dffe_23(pipeline_dffe_23),
	.pipeline_dffe_22(pipeline_dffe_22),
	.pipeline_dffe_21(pipeline_dffe_21),
	.pipeline_dffe_20(pipeline_dffe_20),
	.pipeline_dffe_19(pipeline_dffe_19),
	.pipeline_dffe_18(pipeline_dffe_18),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_11(pipeline_dffe_11),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module nco_test_add_sub_jmh (
	phi_int_arr_reg_31,
	phi_int_arr_reg_30,
	phi_int_arr_reg_29,
	phi_int_arr_reg_28,
	phi_int_arr_reg_27,
	phi_int_arr_reg_26,
	phi_int_arr_reg_25,
	phi_int_arr_reg_24,
	phi_int_arr_reg_23,
	phi_int_arr_reg_22,
	phi_int_arr_reg_21,
	phi_int_arr_reg_20,
	phi_int_arr_reg_19,
	phi_int_arr_reg_18,
	phi_int_arr_reg_17,
	phi_int_arr_reg_16,
	phi_int_arr_reg_15,
	phi_int_arr_reg_14,
	phi_int_arr_reg_13,
	phi_int_arr_reg_12,
	phi_int_arr_reg_11,
	phi_int_arr_reg_10,
	phi_int_arr_reg_9,
	phi_int_arr_reg_8,
	phi_int_arr_reg_7,
	phi_int_arr_reg_6,
	phi_int_arr_reg_5,
	phi_int_arr_reg_4,
	phi_int_arr_reg_3,
	phi_int_arr_reg_2,
	phi_int_arr_reg_1,
	phi_int_arr_reg_0,
	pipeline_dffe_31,
	pipeline_dffe_30,
	pipeline_dffe_29,
	pipeline_dffe_28,
	pipeline_dffe_27,
	pipeline_dffe_26,
	pipeline_dffe_25,
	pipeline_dffe_24,
	pipeline_dffe_23,
	pipeline_dffe_22,
	pipeline_dffe_21,
	pipeline_dffe_20,
	pipeline_dffe_19,
	pipeline_dffe_18,
	pipeline_dffe_17,
	pipeline_dffe_16,
	pipeline_dffe_15,
	pipeline_dffe_14,
	pipeline_dffe_13,
	pipeline_dffe_12,
	pipeline_dffe_11,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	phi_int_arr_reg_31;
input 	phi_int_arr_reg_30;
input 	phi_int_arr_reg_29;
input 	phi_int_arr_reg_28;
input 	phi_int_arr_reg_27;
input 	phi_int_arr_reg_26;
input 	phi_int_arr_reg_25;
input 	phi_int_arr_reg_24;
input 	phi_int_arr_reg_23;
input 	phi_int_arr_reg_22;
input 	phi_int_arr_reg_21;
input 	phi_int_arr_reg_20;
input 	phi_int_arr_reg_19;
input 	phi_int_arr_reg_18;
input 	phi_int_arr_reg_17;
input 	phi_int_arr_reg_16;
input 	phi_int_arr_reg_15;
input 	phi_int_arr_reg_14;
input 	phi_int_arr_reg_13;
input 	phi_int_arr_reg_12;
input 	phi_int_arr_reg_11;
input 	phi_int_arr_reg_10;
input 	phi_int_arr_reg_9;
input 	phi_int_arr_reg_8;
input 	phi_int_arr_reg_7;
input 	phi_int_arr_reg_6;
input 	phi_int_arr_reg_5;
input 	phi_int_arr_reg_4;
input 	phi_int_arr_reg_3;
input 	phi_int_arr_reg_2;
input 	phi_int_arr_reg_1;
input 	phi_int_arr_reg_0;
output 	pipeline_dffe_31;
output 	pipeline_dffe_30;
output 	pipeline_dffe_29;
output 	pipeline_dffe_28;
output 	pipeline_dffe_27;
output 	pipeline_dffe_26;
output 	pipeline_dffe_25;
output 	pipeline_dffe_24;
output 	pipeline_dffe_23;
output 	pipeline_dffe_22;
output 	pipeline_dffe_21;
output 	pipeline_dffe_20;
output 	pipeline_dffe_19;
output 	pipeline_dffe_18;
output 	pipeline_dffe_17;
output 	pipeline_dffe_16;
output 	pipeline_dffe_15;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \op_1~125_sumout ;
wire \pipeline_dffe[0]~q ;
wire \op_1~126 ;
wire \op_1~121_sumout ;
wire \pipeline_dffe[1]~q ;
wire \op_1~122 ;
wire \op_1~117_sumout ;
wire \pipeline_dffe[2]~q ;
wire \op_1~118 ;
wire \op_1~113_sumout ;
wire \pipeline_dffe[3]~q ;
wire \op_1~114 ;
wire \op_1~109_sumout ;
wire \pipeline_dffe[4]~q ;
wire \op_1~110 ;
wire \op_1~105_sumout ;
wire \pipeline_dffe[5]~q ;
wire \op_1~106 ;
wire \op_1~101_sumout ;
wire \pipeline_dffe[6]~q ;
wire \op_1~102 ;
wire \op_1~97_sumout ;
wire \pipeline_dffe[7]~q ;
wire \op_1~98 ;
wire \op_1~93_sumout ;
wire \pipeline_dffe[8]~q ;
wire \op_1~94 ;
wire \op_1~89_sumout ;
wire \pipeline_dffe[9]~q ;
wire \op_1~90 ;
wire \op_1~85_sumout ;
wire \pipeline_dffe[10]~q ;
wire \op_1~86 ;
wire \op_1~82 ;
wire \op_1~78 ;
wire \op_1~74 ;
wire \op_1~70 ;
wire \op_1~66 ;
wire \op_1~62 ;
wire \op_1~58 ;
wire \op_1~54 ;
wire \op_1~50 ;
wire \op_1~46 ;
wire \op_1~42 ;
wire \op_1~38 ;
wire \op_1~34 ;
wire \op_1~30 ;
wire \op_1~26 ;
wire \op_1~22 ;
wire \op_1~18 ;
wire \op_1~14 ;
wire \op_1~10 ;
wire \op_1~6 ;
wire \op_1~1_sumout ;
wire \op_1~5_sumout ;
wire \op_1~9_sumout ;
wire \op_1~13_sumout ;
wire \op_1~17_sumout ;
wire \op_1~21_sumout ;
wire \op_1~25_sumout ;
wire \op_1~29_sumout ;
wire \op_1~33_sumout ;
wire \op_1~37_sumout ;
wire \op_1~41_sumout ;
wire \op_1~45_sumout ;
wire \op_1~49_sumout ;
wire \op_1~53_sumout ;
wire \op_1~57_sumout ;
wire \op_1~61_sumout ;
wire \op_1~65_sumout ;
wire \op_1~69_sumout ;
wire \op_1~73_sumout ;
wire \op_1~77_sumout ;
wire \op_1~81_sumout ;


dffeas \pipeline_dffe[31] (
	.clk(clock),
	.d(\op_1~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_31),
	.prn(vcc));
defparam \pipeline_dffe[31] .is_wysiwyg = "true";
defparam \pipeline_dffe[31] .power_up = "low";

dffeas \pipeline_dffe[30] (
	.clk(clock),
	.d(\op_1~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_30),
	.prn(vcc));
defparam \pipeline_dffe[30] .is_wysiwyg = "true";
defparam \pipeline_dffe[30] .power_up = "low";

dffeas \pipeline_dffe[29] (
	.clk(clock),
	.d(\op_1~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_29),
	.prn(vcc));
defparam \pipeline_dffe[29] .is_wysiwyg = "true";
defparam \pipeline_dffe[29] .power_up = "low";

dffeas \pipeline_dffe[28] (
	.clk(clock),
	.d(\op_1~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_28),
	.prn(vcc));
defparam \pipeline_dffe[28] .is_wysiwyg = "true";
defparam \pipeline_dffe[28] .power_up = "low";

dffeas \pipeline_dffe[27] (
	.clk(clock),
	.d(\op_1~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_27),
	.prn(vcc));
defparam \pipeline_dffe[27] .is_wysiwyg = "true";
defparam \pipeline_dffe[27] .power_up = "low";

dffeas \pipeline_dffe[26] (
	.clk(clock),
	.d(\op_1~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_26),
	.prn(vcc));
defparam \pipeline_dffe[26] .is_wysiwyg = "true";
defparam \pipeline_dffe[26] .power_up = "low";

dffeas \pipeline_dffe[25] (
	.clk(clock),
	.d(\op_1~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_25),
	.prn(vcc));
defparam \pipeline_dffe[25] .is_wysiwyg = "true";
defparam \pipeline_dffe[25] .power_up = "low";

dffeas \pipeline_dffe[24] (
	.clk(clock),
	.d(\op_1~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_24),
	.prn(vcc));
defparam \pipeline_dffe[24] .is_wysiwyg = "true";
defparam \pipeline_dffe[24] .power_up = "low";

dffeas \pipeline_dffe[23] (
	.clk(clock),
	.d(\op_1~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_23),
	.prn(vcc));
defparam \pipeline_dffe[23] .is_wysiwyg = "true";
defparam \pipeline_dffe[23] .power_up = "low";

dffeas \pipeline_dffe[22] (
	.clk(clock),
	.d(\op_1~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_22),
	.prn(vcc));
defparam \pipeline_dffe[22] .is_wysiwyg = "true";
defparam \pipeline_dffe[22] .power_up = "low";

dffeas \pipeline_dffe[21] (
	.clk(clock),
	.d(\op_1~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_21),
	.prn(vcc));
defparam \pipeline_dffe[21] .is_wysiwyg = "true";
defparam \pipeline_dffe[21] .power_up = "low";

dffeas \pipeline_dffe[20] (
	.clk(clock),
	.d(\op_1~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_20),
	.prn(vcc));
defparam \pipeline_dffe[20] .is_wysiwyg = "true";
defparam \pipeline_dffe[20] .power_up = "low";

dffeas \pipeline_dffe[19] (
	.clk(clock),
	.d(\op_1~49_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_19),
	.prn(vcc));
defparam \pipeline_dffe[19] .is_wysiwyg = "true";
defparam \pipeline_dffe[19] .power_up = "low";

dffeas \pipeline_dffe[18] (
	.clk(clock),
	.d(\op_1~53_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_18),
	.prn(vcc));
defparam \pipeline_dffe[18] .is_wysiwyg = "true";
defparam \pipeline_dffe[18] .power_up = "low";

dffeas \pipeline_dffe[17] (
	.clk(clock),
	.d(\op_1~57_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_17),
	.prn(vcc));
defparam \pipeline_dffe[17] .is_wysiwyg = "true";
defparam \pipeline_dffe[17] .power_up = "low";

dffeas \pipeline_dffe[16] (
	.clk(clock),
	.d(\op_1~61_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_16),
	.prn(vcc));
defparam \pipeline_dffe[16] .is_wysiwyg = "true";
defparam \pipeline_dffe[16] .power_up = "low";

dffeas \pipeline_dffe[15] (
	.clk(clock),
	.d(\op_1~65_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_15),
	.prn(vcc));
defparam \pipeline_dffe[15] .is_wysiwyg = "true";
defparam \pipeline_dffe[15] .power_up = "low";

dffeas \pipeline_dffe[14] (
	.clk(clock),
	.d(\op_1~69_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_14),
	.prn(vcc));
defparam \pipeline_dffe[14] .is_wysiwyg = "true";
defparam \pipeline_dffe[14] .power_up = "low";

dffeas \pipeline_dffe[13] (
	.clk(clock),
	.d(\op_1~73_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_13),
	.prn(vcc));
defparam \pipeline_dffe[13] .is_wysiwyg = "true";
defparam \pipeline_dffe[13] .power_up = "low";

dffeas \pipeline_dffe[12] (
	.clk(clock),
	.d(\op_1~77_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_12),
	.prn(vcc));
defparam \pipeline_dffe[12] .is_wysiwyg = "true";
defparam \pipeline_dffe[12] .power_up = "low";

dffeas \pipeline_dffe[11] (
	.clk(clock),
	.d(\op_1~81_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \pipeline_dffe[11] .is_wysiwyg = "true";
defparam \pipeline_dffe[11] .power_up = "low";

arriav_lcell_comb \op_1~125 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_0),
	.datae(gnd),
	.dataf(!\pipeline_dffe[0]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~125_sumout ),
	.cout(\op_1~126 ),
	.shareout());
defparam \op_1~125 .extended_lut = "off";
defparam \op_1~125 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~125 .shared_arith = "off";

dffeas \pipeline_dffe[0] (
	.clk(clock),
	.d(\op_1~125_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[0]~q ),
	.prn(vcc));
defparam \pipeline_dffe[0] .is_wysiwyg = "true";
defparam \pipeline_dffe[0] .power_up = "low";

arriav_lcell_comb \op_1~121 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_1),
	.datae(gnd),
	.dataf(!\pipeline_dffe[1]~q ),
	.datag(gnd),
	.cin(\op_1~126 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~121_sumout ),
	.cout(\op_1~122 ),
	.shareout());
defparam \op_1~121 .extended_lut = "off";
defparam \op_1~121 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~121 .shared_arith = "off";

dffeas \pipeline_dffe[1] (
	.clk(clock),
	.d(\op_1~121_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[1]~q ),
	.prn(vcc));
defparam \pipeline_dffe[1] .is_wysiwyg = "true";
defparam \pipeline_dffe[1] .power_up = "low";

arriav_lcell_comb \op_1~117 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_2),
	.datae(gnd),
	.dataf(!\pipeline_dffe[2]~q ),
	.datag(gnd),
	.cin(\op_1~122 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~117_sumout ),
	.cout(\op_1~118 ),
	.shareout());
defparam \op_1~117 .extended_lut = "off";
defparam \op_1~117 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~117 .shared_arith = "off";

dffeas \pipeline_dffe[2] (
	.clk(clock),
	.d(\op_1~117_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[2]~q ),
	.prn(vcc));
defparam \pipeline_dffe[2] .is_wysiwyg = "true";
defparam \pipeline_dffe[2] .power_up = "low";

arriav_lcell_comb \op_1~113 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_3),
	.datae(gnd),
	.dataf(!\pipeline_dffe[3]~q ),
	.datag(gnd),
	.cin(\op_1~118 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~113_sumout ),
	.cout(\op_1~114 ),
	.shareout());
defparam \op_1~113 .extended_lut = "off";
defparam \op_1~113 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~113 .shared_arith = "off";

dffeas \pipeline_dffe[3] (
	.clk(clock),
	.d(\op_1~113_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[3]~q ),
	.prn(vcc));
defparam \pipeline_dffe[3] .is_wysiwyg = "true";
defparam \pipeline_dffe[3] .power_up = "low";

arriav_lcell_comb \op_1~109 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_4),
	.datae(gnd),
	.dataf(!\pipeline_dffe[4]~q ),
	.datag(gnd),
	.cin(\op_1~114 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~109_sumout ),
	.cout(\op_1~110 ),
	.shareout());
defparam \op_1~109 .extended_lut = "off";
defparam \op_1~109 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~109 .shared_arith = "off";

dffeas \pipeline_dffe[4] (
	.clk(clock),
	.d(\op_1~109_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[4]~q ),
	.prn(vcc));
defparam \pipeline_dffe[4] .is_wysiwyg = "true";
defparam \pipeline_dffe[4] .power_up = "low";

arriav_lcell_comb \op_1~105 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_5),
	.datae(gnd),
	.dataf(!\pipeline_dffe[5]~q ),
	.datag(gnd),
	.cin(\op_1~110 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~105_sumout ),
	.cout(\op_1~106 ),
	.shareout());
defparam \op_1~105 .extended_lut = "off";
defparam \op_1~105 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~105 .shared_arith = "off";

dffeas \pipeline_dffe[5] (
	.clk(clock),
	.d(\op_1~105_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[5]~q ),
	.prn(vcc));
defparam \pipeline_dffe[5] .is_wysiwyg = "true";
defparam \pipeline_dffe[5] .power_up = "low";

arriav_lcell_comb \op_1~101 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_6),
	.datae(gnd),
	.dataf(!\pipeline_dffe[6]~q ),
	.datag(gnd),
	.cin(\op_1~106 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~101_sumout ),
	.cout(\op_1~102 ),
	.shareout());
defparam \op_1~101 .extended_lut = "off";
defparam \op_1~101 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~101 .shared_arith = "off";

dffeas \pipeline_dffe[6] (
	.clk(clock),
	.d(\op_1~101_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[6]~q ),
	.prn(vcc));
defparam \pipeline_dffe[6] .is_wysiwyg = "true";
defparam \pipeline_dffe[6] .power_up = "low";

arriav_lcell_comb \op_1~97 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_7),
	.datae(gnd),
	.dataf(!\pipeline_dffe[7]~q ),
	.datag(gnd),
	.cin(\op_1~102 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~97_sumout ),
	.cout(\op_1~98 ),
	.shareout());
defparam \op_1~97 .extended_lut = "off";
defparam \op_1~97 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~97 .shared_arith = "off";

dffeas \pipeline_dffe[7] (
	.clk(clock),
	.d(\op_1~97_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[7]~q ),
	.prn(vcc));
defparam \pipeline_dffe[7] .is_wysiwyg = "true";
defparam \pipeline_dffe[7] .power_up = "low";

arriav_lcell_comb \op_1~93 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_8),
	.datae(gnd),
	.dataf(!\pipeline_dffe[8]~q ),
	.datag(gnd),
	.cin(\op_1~98 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~93_sumout ),
	.cout(\op_1~94 ),
	.shareout());
defparam \op_1~93 .extended_lut = "off";
defparam \op_1~93 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~93 .shared_arith = "off";

dffeas \pipeline_dffe[8] (
	.clk(clock),
	.d(\op_1~93_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[8]~q ),
	.prn(vcc));
defparam \pipeline_dffe[8] .is_wysiwyg = "true";
defparam \pipeline_dffe[8] .power_up = "low";

arriav_lcell_comb \op_1~89 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_9),
	.datae(gnd),
	.dataf(!\pipeline_dffe[9]~q ),
	.datag(gnd),
	.cin(\op_1~94 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~89_sumout ),
	.cout(\op_1~90 ),
	.shareout());
defparam \op_1~89 .extended_lut = "off";
defparam \op_1~89 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~89 .shared_arith = "off";

dffeas \pipeline_dffe[9] (
	.clk(clock),
	.d(\op_1~89_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[9]~q ),
	.prn(vcc));
defparam \pipeline_dffe[9] .is_wysiwyg = "true";
defparam \pipeline_dffe[9] .power_up = "low";

arriav_lcell_comb \op_1~85 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_10),
	.datae(gnd),
	.dataf(!\pipeline_dffe[10]~q ),
	.datag(gnd),
	.cin(\op_1~90 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~85_sumout ),
	.cout(\op_1~86 ),
	.shareout());
defparam \op_1~85 .extended_lut = "off";
defparam \op_1~85 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~85 .shared_arith = "off";

dffeas \pipeline_dffe[10] (
	.clk(clock),
	.d(\op_1~85_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(\pipeline_dffe[10]~q ),
	.prn(vcc));
defparam \pipeline_dffe[10] .is_wysiwyg = "true";
defparam \pipeline_dffe[10] .power_up = "low";

arriav_lcell_comb \op_1~81 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_11),
	.datae(gnd),
	.dataf(!pipeline_dffe_11),
	.datag(gnd),
	.cin(\op_1~86 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~81_sumout ),
	.cout(\op_1~82 ),
	.shareout());
defparam \op_1~81 .extended_lut = "off";
defparam \op_1~81 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~81 .shared_arith = "off";

arriav_lcell_comb \op_1~77 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_12),
	.datae(gnd),
	.dataf(!pipeline_dffe_12),
	.datag(gnd),
	.cin(\op_1~82 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~77_sumout ),
	.cout(\op_1~78 ),
	.shareout());
defparam \op_1~77 .extended_lut = "off";
defparam \op_1~77 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~77 .shared_arith = "off";

arriav_lcell_comb \op_1~73 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_13),
	.datae(gnd),
	.dataf(!pipeline_dffe_13),
	.datag(gnd),
	.cin(\op_1~78 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~73_sumout ),
	.cout(\op_1~74 ),
	.shareout());
defparam \op_1~73 .extended_lut = "off";
defparam \op_1~73 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~73 .shared_arith = "off";

arriav_lcell_comb \op_1~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_14),
	.datae(gnd),
	.dataf(!pipeline_dffe_14),
	.datag(gnd),
	.cin(\op_1~74 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~69_sumout ),
	.cout(\op_1~70 ),
	.shareout());
defparam \op_1~69 .extended_lut = "off";
defparam \op_1~69 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~69 .shared_arith = "off";

arriav_lcell_comb \op_1~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_15),
	.datae(gnd),
	.dataf(!pipeline_dffe_15),
	.datag(gnd),
	.cin(\op_1~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~65_sumout ),
	.cout(\op_1~66 ),
	.shareout());
defparam \op_1~65 .extended_lut = "off";
defparam \op_1~65 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~65 .shared_arith = "off";

arriav_lcell_comb \op_1~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_16),
	.datae(gnd),
	.dataf(!pipeline_dffe_16),
	.datag(gnd),
	.cin(\op_1~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~61_sumout ),
	.cout(\op_1~62 ),
	.shareout());
defparam \op_1~61 .extended_lut = "off";
defparam \op_1~61 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~61 .shared_arith = "off";

arriav_lcell_comb \op_1~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_17),
	.datae(gnd),
	.dataf(!pipeline_dffe_17),
	.datag(gnd),
	.cin(\op_1~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~57_sumout ),
	.cout(\op_1~58 ),
	.shareout());
defparam \op_1~57 .extended_lut = "off";
defparam \op_1~57 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~57 .shared_arith = "off";

arriav_lcell_comb \op_1~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_18),
	.datae(gnd),
	.dataf(!pipeline_dffe_18),
	.datag(gnd),
	.cin(\op_1~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~53_sumout ),
	.cout(\op_1~54 ),
	.shareout());
defparam \op_1~53 .extended_lut = "off";
defparam \op_1~53 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~53 .shared_arith = "off";

arriav_lcell_comb \op_1~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_19),
	.datae(gnd),
	.dataf(!pipeline_dffe_19),
	.datag(gnd),
	.cin(\op_1~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~49_sumout ),
	.cout(\op_1~50 ),
	.shareout());
defparam \op_1~49 .extended_lut = "off";
defparam \op_1~49 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~49 .shared_arith = "off";

arriav_lcell_comb \op_1~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_20),
	.datae(gnd),
	.dataf(!pipeline_dffe_20),
	.datag(gnd),
	.cin(\op_1~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~45_sumout ),
	.cout(\op_1~46 ),
	.shareout());
defparam \op_1~45 .extended_lut = "off";
defparam \op_1~45 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~45 .shared_arith = "off";

arriav_lcell_comb \op_1~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_21),
	.datae(gnd),
	.dataf(!pipeline_dffe_21),
	.datag(gnd),
	.cin(\op_1~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~41_sumout ),
	.cout(\op_1~42 ),
	.shareout());
defparam \op_1~41 .extended_lut = "off";
defparam \op_1~41 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~41 .shared_arith = "off";

arriav_lcell_comb \op_1~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_22),
	.datae(gnd),
	.dataf(!pipeline_dffe_22),
	.datag(gnd),
	.cin(\op_1~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~37_sumout ),
	.cout(\op_1~38 ),
	.shareout());
defparam \op_1~37 .extended_lut = "off";
defparam \op_1~37 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~37 .shared_arith = "off";

arriav_lcell_comb \op_1~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_23),
	.datae(gnd),
	.dataf(!pipeline_dffe_23),
	.datag(gnd),
	.cin(\op_1~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~33_sumout ),
	.cout(\op_1~34 ),
	.shareout());
defparam \op_1~33 .extended_lut = "off";
defparam \op_1~33 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~33 .shared_arith = "off";

arriav_lcell_comb \op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_24),
	.datae(gnd),
	.dataf(!pipeline_dffe_24),
	.datag(gnd),
	.cin(\op_1~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~29_sumout ),
	.cout(\op_1~30 ),
	.shareout());
defparam \op_1~29 .extended_lut = "off";
defparam \op_1~29 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~29 .shared_arith = "off";

arriav_lcell_comb \op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_25),
	.datae(gnd),
	.dataf(!pipeline_dffe_25),
	.datag(gnd),
	.cin(\op_1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~25_sumout ),
	.cout(\op_1~26 ),
	.shareout());
defparam \op_1~25 .extended_lut = "off";
defparam \op_1~25 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~25 .shared_arith = "off";

arriav_lcell_comb \op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_26),
	.datae(gnd),
	.dataf(!pipeline_dffe_26),
	.datag(gnd),
	.cin(\op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~21_sumout ),
	.cout(\op_1~22 ),
	.shareout());
defparam \op_1~21 .extended_lut = "off";
defparam \op_1~21 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~21 .shared_arith = "off";

arriav_lcell_comb \op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_27),
	.datae(gnd),
	.dataf(!pipeline_dffe_27),
	.datag(gnd),
	.cin(\op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~17_sumout ),
	.cout(\op_1~18 ),
	.shareout());
defparam \op_1~17 .extended_lut = "off";
defparam \op_1~17 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~17 .shared_arith = "off";

arriav_lcell_comb \op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_28),
	.datae(gnd),
	.dataf(!pipeline_dffe_28),
	.datag(gnd),
	.cin(\op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~13_sumout ),
	.cout(\op_1~14 ),
	.shareout());
defparam \op_1~13 .extended_lut = "off";
defparam \op_1~13 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~13 .shared_arith = "off";

arriav_lcell_comb \op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_29),
	.datae(gnd),
	.dataf(!pipeline_dffe_29),
	.datag(gnd),
	.cin(\op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~9_sumout ),
	.cout(\op_1~10 ),
	.shareout());
defparam \op_1~9 .extended_lut = "off";
defparam \op_1~9 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~9 .shared_arith = "off";

arriav_lcell_comb \op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_30),
	.datae(gnd),
	.dataf(!pipeline_dffe_30),
	.datag(gnd),
	.cin(\op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~5_sumout ),
	.cout(\op_1~6 ),
	.shareout());
defparam \op_1~5 .extended_lut = "off";
defparam \op_1~5 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~5 .shared_arith = "off";

arriav_lcell_comb \op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!phi_int_arr_reg_31),
	.datae(gnd),
	.dataf(!pipeline_dffe_31),
	.datag(gnd),
	.cin(\op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~1_sumout ),
	.cout(),
	.shareout());
defparam \op_1~1 .extended_lut = "off";
defparam \op_1~1 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~1 .shared_arith = "off";

endmodule

module nco_test_asj_crd_par (
	sin_o_0,
	sin_o_1,
	sin_o_2,
	sin_o_3,
	sin_o_4,
	sin_o_5,
	sin_o_6,
	sin_o_7,
	sin_o_8,
	sin_o_9,
	sin_o_10,
	sin_o_11,
	sin_o_12,
	sin_o_13,
	sin_o_14,
	sin_o_15,
	sin_o_16,
	sin_o_17,
	cos_o_0,
	cos_o_1,
	cos_o_2,
	cos_o_3,
	cos_o_4,
	cos_o_5,
	cos_o_6,
	cos_o_7,
	cos_o_8,
	cos_o_9,
	cos_o_10,
	cos_o_11,
	cos_o_12,
	cos_o_13,
	cos_o_14,
	cos_o_15,
	cos_o_16,
	cos_o_17,
	cordic_y_res_d_0,
	cordic_y_res_2c_0,
	cordic_x_res_d_0,
	cordic_x_res_2c_0,
	seg_rot_1,
	seg_rot_0,
	cordic_y_res_d_1,
	cordic_y_res_2c_1,
	cordic_x_res_d_1,
	cordic_x_res_2c_1,
	cordic_y_res_d_2,
	cordic_y_res_2c_2,
	cordic_x_res_d_2,
	cordic_x_res_2c_2,
	cordic_y_res_d_3,
	cordic_y_res_2c_3,
	cordic_x_res_d_3,
	cordic_x_res_2c_3,
	cordic_y_res_d_4,
	cordic_y_res_2c_4,
	cordic_x_res_d_4,
	cordic_x_res_2c_4,
	cordic_y_res_d_5,
	cordic_y_res_2c_5,
	cordic_x_res_d_5,
	cordic_x_res_2c_5,
	cordic_y_res_d_6,
	cordic_y_res_2c_6,
	cordic_x_res_d_6,
	cordic_x_res_2c_6,
	cordic_y_res_d_7,
	cordic_y_res_2c_7,
	cordic_x_res_d_7,
	cordic_x_res_2c_7,
	cordic_y_res_d_8,
	cordic_y_res_2c_8,
	cordic_x_res_d_8,
	cordic_x_res_2c_8,
	cordic_y_res_d_9,
	cordic_y_res_2c_9,
	cordic_x_res_d_9,
	cordic_x_res_2c_9,
	cordic_y_res_d_10,
	cordic_y_res_2c_10,
	cordic_x_res_d_10,
	cordic_x_res_2c_10,
	cordic_y_res_d_11,
	cordic_y_res_2c_11,
	cordic_x_res_d_11,
	cordic_x_res_2c_11,
	cordic_y_res_d_12,
	cordic_y_res_2c_12,
	cordic_x_res_d_12,
	cordic_x_res_2c_12,
	cordic_y_res_d_13,
	cordic_y_res_2c_13,
	cordic_x_res_d_13,
	cordic_x_res_2c_13,
	cordic_y_res_d_14,
	cordic_y_res_2c_14,
	cordic_x_res_d_14,
	cordic_x_res_2c_14,
	cordic_y_res_d_15,
	cordic_y_res_2c_15,
	cordic_x_res_d_15,
	cordic_x_res_2c_15,
	cordic_y_res_d_16,
	cordic_y_res_2c_16,
	cordic_x_res_d_16,
	cordic_x_res_2c_16,
	cordic_y_res_d_17,
	cordic_y_res_2c_17,
	cordic_x_res_d_17,
	cordic_x_res_2c_17,
	sin_o_01,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	sin_o_0;
output 	sin_o_1;
output 	sin_o_2;
output 	sin_o_3;
output 	sin_o_4;
output 	sin_o_5;
output 	sin_o_6;
output 	sin_o_7;
output 	sin_o_8;
output 	sin_o_9;
output 	sin_o_10;
output 	sin_o_11;
output 	sin_o_12;
output 	sin_o_13;
output 	sin_o_14;
output 	sin_o_15;
output 	sin_o_16;
output 	sin_o_17;
output 	cos_o_0;
output 	cos_o_1;
output 	cos_o_2;
output 	cos_o_3;
output 	cos_o_4;
output 	cos_o_5;
output 	cos_o_6;
output 	cos_o_7;
output 	cos_o_8;
output 	cos_o_9;
output 	cos_o_10;
output 	cos_o_11;
output 	cos_o_12;
output 	cos_o_13;
output 	cos_o_14;
output 	cos_o_15;
output 	cos_o_16;
output 	cos_o_17;
input 	cordic_y_res_d_0;
input 	cordic_y_res_2c_0;
input 	cordic_x_res_d_0;
input 	cordic_x_res_2c_0;
input 	seg_rot_1;
input 	seg_rot_0;
input 	cordic_y_res_d_1;
input 	cordic_y_res_2c_1;
input 	cordic_x_res_d_1;
input 	cordic_x_res_2c_1;
input 	cordic_y_res_d_2;
input 	cordic_y_res_2c_2;
input 	cordic_x_res_d_2;
input 	cordic_x_res_2c_2;
input 	cordic_y_res_d_3;
input 	cordic_y_res_2c_3;
input 	cordic_x_res_d_3;
input 	cordic_x_res_2c_3;
input 	cordic_y_res_d_4;
input 	cordic_y_res_2c_4;
input 	cordic_x_res_d_4;
input 	cordic_x_res_2c_4;
input 	cordic_y_res_d_5;
input 	cordic_y_res_2c_5;
input 	cordic_x_res_d_5;
input 	cordic_x_res_2c_5;
input 	cordic_y_res_d_6;
input 	cordic_y_res_2c_6;
input 	cordic_x_res_d_6;
input 	cordic_x_res_2c_6;
input 	cordic_y_res_d_7;
input 	cordic_y_res_2c_7;
input 	cordic_x_res_d_7;
input 	cordic_x_res_2c_7;
input 	cordic_y_res_d_8;
input 	cordic_y_res_2c_8;
input 	cordic_x_res_d_8;
input 	cordic_x_res_2c_8;
input 	cordic_y_res_d_9;
input 	cordic_y_res_2c_9;
input 	cordic_x_res_d_9;
input 	cordic_x_res_2c_9;
input 	cordic_y_res_d_10;
input 	cordic_y_res_2c_10;
input 	cordic_x_res_d_10;
input 	cordic_x_res_2c_10;
input 	cordic_y_res_d_11;
input 	cordic_y_res_2c_11;
input 	cordic_x_res_d_11;
input 	cordic_x_res_2c_11;
input 	cordic_y_res_d_12;
input 	cordic_y_res_2c_12;
input 	cordic_x_res_d_12;
input 	cordic_x_res_2c_12;
input 	cordic_y_res_d_13;
input 	cordic_y_res_2c_13;
input 	cordic_x_res_d_13;
input 	cordic_x_res_2c_13;
input 	cordic_y_res_d_14;
input 	cordic_y_res_2c_14;
input 	cordic_x_res_d_14;
input 	cordic_x_res_2c_14;
input 	cordic_y_res_d_15;
input 	cordic_y_res_2c_15;
input 	cordic_x_res_d_15;
input 	cordic_x_res_2c_15;
input 	cordic_y_res_d_16;
input 	cordic_y_res_2c_16;
input 	cordic_x_res_d_16;
input 	cordic_x_res_2c_16;
input 	cordic_y_res_d_17;
input 	cordic_y_res_2c_17;
input 	cordic_x_res_d_17;
input 	cordic_x_res_2c_17;
input 	sin_o_01;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \sin_o~0_combout ;
wire \sin_o~1_combout ;
wire \sin_o~2_combout ;
wire \sin_o~3_combout ;
wire \sin_o~4_combout ;
wire \sin_o~5_combout ;
wire \sin_o~6_combout ;
wire \sin_o~7_combout ;
wire \sin_o~8_combout ;
wire \sin_o~9_combout ;
wire \sin_o~10_combout ;
wire \sin_o~11_combout ;
wire \sin_o~12_combout ;
wire \sin_o~13_combout ;
wire \sin_o~14_combout ;
wire \sin_o~15_combout ;
wire \sin_o~16_combout ;
wire \sin_o~17_combout ;
wire \cos_o~0_combout ;
wire \cos_o~1_combout ;
wire \cos_o~2_combout ;
wire \cos_o~3_combout ;
wire \cos_o~4_combout ;
wire \cos_o~5_combout ;
wire \cos_o~6_combout ;
wire \cos_o~7_combout ;
wire \cos_o~8_combout ;
wire \cos_o~9_combout ;
wire \cos_o~10_combout ;
wire \cos_o~11_combout ;
wire \cos_o~12_combout ;
wire \cos_o~13_combout ;
wire \cos_o~14_combout ;
wire \cos_o~15_combout ;
wire \cos_o~16_combout ;
wire \cos_o~17_combout ;


dffeas \sin_o[0] (
	.clk(clk),
	.d(\sin_o~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_01),
	.q(sin_o_0),
	.prn(vcc));
defparam \sin_o[0] .is_wysiwyg = "true";
defparam \sin_o[0] .power_up = "low";

dffeas \sin_o[1] (
	.clk(clk),
	.d(\sin_o~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_01),
	.q(sin_o_1),
	.prn(vcc));
defparam \sin_o[1] .is_wysiwyg = "true";
defparam \sin_o[1] .power_up = "low";

dffeas \sin_o[2] (
	.clk(clk),
	.d(\sin_o~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_01),
	.q(sin_o_2),
	.prn(vcc));
defparam \sin_o[2] .is_wysiwyg = "true";
defparam \sin_o[2] .power_up = "low";

dffeas \sin_o[3] (
	.clk(clk),
	.d(\sin_o~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_01),
	.q(sin_o_3),
	.prn(vcc));
defparam \sin_o[3] .is_wysiwyg = "true";
defparam \sin_o[3] .power_up = "low";

dffeas \sin_o[4] (
	.clk(clk),
	.d(\sin_o~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_01),
	.q(sin_o_4),
	.prn(vcc));
defparam \sin_o[4] .is_wysiwyg = "true";
defparam \sin_o[4] .power_up = "low";

dffeas \sin_o[5] (
	.clk(clk),
	.d(\sin_o~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_01),
	.q(sin_o_5),
	.prn(vcc));
defparam \sin_o[5] .is_wysiwyg = "true";
defparam \sin_o[5] .power_up = "low";

dffeas \sin_o[6] (
	.clk(clk),
	.d(\sin_o~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_01),
	.q(sin_o_6),
	.prn(vcc));
defparam \sin_o[6] .is_wysiwyg = "true";
defparam \sin_o[6] .power_up = "low";

dffeas \sin_o[7] (
	.clk(clk),
	.d(\sin_o~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_01),
	.q(sin_o_7),
	.prn(vcc));
defparam \sin_o[7] .is_wysiwyg = "true";
defparam \sin_o[7] .power_up = "low";

dffeas \sin_o[8] (
	.clk(clk),
	.d(\sin_o~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_01),
	.q(sin_o_8),
	.prn(vcc));
defparam \sin_o[8] .is_wysiwyg = "true";
defparam \sin_o[8] .power_up = "low";

dffeas \sin_o[9] (
	.clk(clk),
	.d(\sin_o~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_01),
	.q(sin_o_9),
	.prn(vcc));
defparam \sin_o[9] .is_wysiwyg = "true";
defparam \sin_o[9] .power_up = "low";

dffeas \sin_o[10] (
	.clk(clk),
	.d(\sin_o~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_01),
	.q(sin_o_10),
	.prn(vcc));
defparam \sin_o[10] .is_wysiwyg = "true";
defparam \sin_o[10] .power_up = "low";

dffeas \sin_o[11] (
	.clk(clk),
	.d(\sin_o~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_01),
	.q(sin_o_11),
	.prn(vcc));
defparam \sin_o[11] .is_wysiwyg = "true";
defparam \sin_o[11] .power_up = "low";

dffeas \sin_o[12] (
	.clk(clk),
	.d(\sin_o~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_01),
	.q(sin_o_12),
	.prn(vcc));
defparam \sin_o[12] .is_wysiwyg = "true";
defparam \sin_o[12] .power_up = "low";

dffeas \sin_o[13] (
	.clk(clk),
	.d(\sin_o~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_01),
	.q(sin_o_13),
	.prn(vcc));
defparam \sin_o[13] .is_wysiwyg = "true";
defparam \sin_o[13] .power_up = "low";

dffeas \sin_o[14] (
	.clk(clk),
	.d(\sin_o~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_01),
	.q(sin_o_14),
	.prn(vcc));
defparam \sin_o[14] .is_wysiwyg = "true";
defparam \sin_o[14] .power_up = "low";

dffeas \sin_o[15] (
	.clk(clk),
	.d(\sin_o~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_01),
	.q(sin_o_15),
	.prn(vcc));
defparam \sin_o[15] .is_wysiwyg = "true";
defparam \sin_o[15] .power_up = "low";

dffeas \sin_o[16] (
	.clk(clk),
	.d(\sin_o~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_01),
	.q(sin_o_16),
	.prn(vcc));
defparam \sin_o[16] .is_wysiwyg = "true";
defparam \sin_o[16] .power_up = "low";

dffeas \sin_o[17] (
	.clk(clk),
	.d(\sin_o~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_01),
	.q(sin_o_17),
	.prn(vcc));
defparam \sin_o[17] .is_wysiwyg = "true";
defparam \sin_o[17] .power_up = "low";

dffeas \cos_o[0] (
	.clk(clk),
	.d(\cos_o~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_01),
	.q(cos_o_0),
	.prn(vcc));
defparam \cos_o[0] .is_wysiwyg = "true";
defparam \cos_o[0] .power_up = "low";

dffeas \cos_o[1] (
	.clk(clk),
	.d(\cos_o~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_01),
	.q(cos_o_1),
	.prn(vcc));
defparam \cos_o[1] .is_wysiwyg = "true";
defparam \cos_o[1] .power_up = "low";

dffeas \cos_o[2] (
	.clk(clk),
	.d(\cos_o~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_01),
	.q(cos_o_2),
	.prn(vcc));
defparam \cos_o[2] .is_wysiwyg = "true";
defparam \cos_o[2] .power_up = "low";

dffeas \cos_o[3] (
	.clk(clk),
	.d(\cos_o~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_01),
	.q(cos_o_3),
	.prn(vcc));
defparam \cos_o[3] .is_wysiwyg = "true";
defparam \cos_o[3] .power_up = "low";

dffeas \cos_o[4] (
	.clk(clk),
	.d(\cos_o~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_01),
	.q(cos_o_4),
	.prn(vcc));
defparam \cos_o[4] .is_wysiwyg = "true";
defparam \cos_o[4] .power_up = "low";

dffeas \cos_o[5] (
	.clk(clk),
	.d(\cos_o~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_01),
	.q(cos_o_5),
	.prn(vcc));
defparam \cos_o[5] .is_wysiwyg = "true";
defparam \cos_o[5] .power_up = "low";

dffeas \cos_o[6] (
	.clk(clk),
	.d(\cos_o~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_01),
	.q(cos_o_6),
	.prn(vcc));
defparam \cos_o[6] .is_wysiwyg = "true";
defparam \cos_o[6] .power_up = "low";

dffeas \cos_o[7] (
	.clk(clk),
	.d(\cos_o~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_01),
	.q(cos_o_7),
	.prn(vcc));
defparam \cos_o[7] .is_wysiwyg = "true";
defparam \cos_o[7] .power_up = "low";

dffeas \cos_o[8] (
	.clk(clk),
	.d(\cos_o~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_01),
	.q(cos_o_8),
	.prn(vcc));
defparam \cos_o[8] .is_wysiwyg = "true";
defparam \cos_o[8] .power_up = "low";

dffeas \cos_o[9] (
	.clk(clk),
	.d(\cos_o~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_01),
	.q(cos_o_9),
	.prn(vcc));
defparam \cos_o[9] .is_wysiwyg = "true";
defparam \cos_o[9] .power_up = "low";

dffeas \cos_o[10] (
	.clk(clk),
	.d(\cos_o~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_01),
	.q(cos_o_10),
	.prn(vcc));
defparam \cos_o[10] .is_wysiwyg = "true";
defparam \cos_o[10] .power_up = "low";

dffeas \cos_o[11] (
	.clk(clk),
	.d(\cos_o~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_01),
	.q(cos_o_11),
	.prn(vcc));
defparam \cos_o[11] .is_wysiwyg = "true";
defparam \cos_o[11] .power_up = "low";

dffeas \cos_o[12] (
	.clk(clk),
	.d(\cos_o~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_01),
	.q(cos_o_12),
	.prn(vcc));
defparam \cos_o[12] .is_wysiwyg = "true";
defparam \cos_o[12] .power_up = "low";

dffeas \cos_o[13] (
	.clk(clk),
	.d(\cos_o~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_01),
	.q(cos_o_13),
	.prn(vcc));
defparam \cos_o[13] .is_wysiwyg = "true";
defparam \cos_o[13] .power_up = "low";

dffeas \cos_o[14] (
	.clk(clk),
	.d(\cos_o~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_01),
	.q(cos_o_14),
	.prn(vcc));
defparam \cos_o[14] .is_wysiwyg = "true";
defparam \cos_o[14] .power_up = "low";

dffeas \cos_o[15] (
	.clk(clk),
	.d(\cos_o~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_01),
	.q(cos_o_15),
	.prn(vcc));
defparam \cos_o[15] .is_wysiwyg = "true";
defparam \cos_o[15] .power_up = "low";

dffeas \cos_o[16] (
	.clk(clk),
	.d(\cos_o~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_01),
	.q(cos_o_16),
	.prn(vcc));
defparam \cos_o[16] .is_wysiwyg = "true";
defparam \cos_o[16] .power_up = "low";

dffeas \cos_o[17] (
	.clk(clk),
	.d(\cos_o~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_01),
	.q(cos_o_17),
	.prn(vcc));
defparam \cos_o[17] .is_wysiwyg = "true";
defparam \cos_o[17] .power_up = "low";

arriav_lcell_comb \sin_o~0 (
	.dataa(!cordic_y_res_d_0),
	.datab(!cordic_y_res_2c_0),
	.datac(!cordic_x_res_d_0),
	.datad(!cordic_x_res_2c_0),
	.datae(!seg_rot_1),
	.dataf(!seg_rot_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sin_o~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sin_o~0 .extended_lut = "off";
defparam \sin_o~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \sin_o~0 .shared_arith = "off";

arriav_lcell_comb \sin_o~1 (
	.dataa(!cordic_y_res_d_1),
	.datab(!cordic_y_res_2c_1),
	.datac(!cordic_x_res_d_1),
	.datad(!cordic_x_res_2c_1),
	.datae(!seg_rot_1),
	.dataf(!seg_rot_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sin_o~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sin_o~1 .extended_lut = "off";
defparam \sin_o~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \sin_o~1 .shared_arith = "off";

arriav_lcell_comb \sin_o~2 (
	.dataa(!cordic_y_res_d_2),
	.datab(!cordic_y_res_2c_2),
	.datac(!cordic_x_res_d_2),
	.datad(!cordic_x_res_2c_2),
	.datae(!seg_rot_1),
	.dataf(!seg_rot_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sin_o~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sin_o~2 .extended_lut = "off";
defparam \sin_o~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \sin_o~2 .shared_arith = "off";

arriav_lcell_comb \sin_o~3 (
	.dataa(!cordic_y_res_d_3),
	.datab(!cordic_y_res_2c_3),
	.datac(!cordic_x_res_d_3),
	.datad(!cordic_x_res_2c_3),
	.datae(!seg_rot_1),
	.dataf(!seg_rot_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sin_o~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sin_o~3 .extended_lut = "off";
defparam \sin_o~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \sin_o~3 .shared_arith = "off";

arriav_lcell_comb \sin_o~4 (
	.dataa(!cordic_y_res_d_4),
	.datab(!cordic_y_res_2c_4),
	.datac(!cordic_x_res_d_4),
	.datad(!cordic_x_res_2c_4),
	.datae(!seg_rot_1),
	.dataf(!seg_rot_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sin_o~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sin_o~4 .extended_lut = "off";
defparam \sin_o~4 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \sin_o~4 .shared_arith = "off";

arriav_lcell_comb \sin_o~5 (
	.dataa(!cordic_y_res_d_5),
	.datab(!cordic_y_res_2c_5),
	.datac(!cordic_x_res_d_5),
	.datad(!cordic_x_res_2c_5),
	.datae(!seg_rot_1),
	.dataf(!seg_rot_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sin_o~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sin_o~5 .extended_lut = "off";
defparam \sin_o~5 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \sin_o~5 .shared_arith = "off";

arriav_lcell_comb \sin_o~6 (
	.dataa(!cordic_y_res_d_6),
	.datab(!cordic_y_res_2c_6),
	.datac(!cordic_x_res_d_6),
	.datad(!cordic_x_res_2c_6),
	.datae(!seg_rot_1),
	.dataf(!seg_rot_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sin_o~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sin_o~6 .extended_lut = "off";
defparam \sin_o~6 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \sin_o~6 .shared_arith = "off";

arriav_lcell_comb \sin_o~7 (
	.dataa(!cordic_y_res_d_7),
	.datab(!cordic_y_res_2c_7),
	.datac(!cordic_x_res_d_7),
	.datad(!cordic_x_res_2c_7),
	.datae(!seg_rot_1),
	.dataf(!seg_rot_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sin_o~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sin_o~7 .extended_lut = "off";
defparam \sin_o~7 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \sin_o~7 .shared_arith = "off";

arriav_lcell_comb \sin_o~8 (
	.dataa(!cordic_y_res_d_8),
	.datab(!cordic_y_res_2c_8),
	.datac(!cordic_x_res_d_8),
	.datad(!cordic_x_res_2c_8),
	.datae(!seg_rot_1),
	.dataf(!seg_rot_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sin_o~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sin_o~8 .extended_lut = "off";
defparam \sin_o~8 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \sin_o~8 .shared_arith = "off";

arriav_lcell_comb \sin_o~9 (
	.dataa(!cordic_y_res_d_9),
	.datab(!cordic_y_res_2c_9),
	.datac(!cordic_x_res_d_9),
	.datad(!cordic_x_res_2c_9),
	.datae(!seg_rot_1),
	.dataf(!seg_rot_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sin_o~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sin_o~9 .extended_lut = "off";
defparam \sin_o~9 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \sin_o~9 .shared_arith = "off";

arriav_lcell_comb \sin_o~10 (
	.dataa(!cordic_y_res_d_10),
	.datab(!cordic_y_res_2c_10),
	.datac(!cordic_x_res_d_10),
	.datad(!cordic_x_res_2c_10),
	.datae(!seg_rot_1),
	.dataf(!seg_rot_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sin_o~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sin_o~10 .extended_lut = "off";
defparam \sin_o~10 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \sin_o~10 .shared_arith = "off";

arriav_lcell_comb \sin_o~11 (
	.dataa(!cordic_y_res_d_11),
	.datab(!cordic_y_res_2c_11),
	.datac(!cordic_x_res_d_11),
	.datad(!cordic_x_res_2c_11),
	.datae(!seg_rot_1),
	.dataf(!seg_rot_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sin_o~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sin_o~11 .extended_lut = "off";
defparam \sin_o~11 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \sin_o~11 .shared_arith = "off";

arriav_lcell_comb \sin_o~12 (
	.dataa(!cordic_y_res_d_12),
	.datab(!cordic_y_res_2c_12),
	.datac(!cordic_x_res_d_12),
	.datad(!cordic_x_res_2c_12),
	.datae(!seg_rot_1),
	.dataf(!seg_rot_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sin_o~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sin_o~12 .extended_lut = "off";
defparam \sin_o~12 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \sin_o~12 .shared_arith = "off";

arriav_lcell_comb \sin_o~13 (
	.dataa(!cordic_y_res_d_13),
	.datab(!cordic_y_res_2c_13),
	.datac(!cordic_x_res_d_13),
	.datad(!cordic_x_res_2c_13),
	.datae(!seg_rot_1),
	.dataf(!seg_rot_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sin_o~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sin_o~13 .extended_lut = "off";
defparam \sin_o~13 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \sin_o~13 .shared_arith = "off";

arriav_lcell_comb \sin_o~14 (
	.dataa(!cordic_y_res_d_14),
	.datab(!cordic_y_res_2c_14),
	.datac(!cordic_x_res_d_14),
	.datad(!cordic_x_res_2c_14),
	.datae(!seg_rot_1),
	.dataf(!seg_rot_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sin_o~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sin_o~14 .extended_lut = "off";
defparam \sin_o~14 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \sin_o~14 .shared_arith = "off";

arriav_lcell_comb \sin_o~15 (
	.dataa(!cordic_y_res_d_15),
	.datab(!cordic_y_res_2c_15),
	.datac(!cordic_x_res_d_15),
	.datad(!cordic_x_res_2c_15),
	.datae(!seg_rot_1),
	.dataf(!seg_rot_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sin_o~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sin_o~15 .extended_lut = "off";
defparam \sin_o~15 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \sin_o~15 .shared_arith = "off";

arriav_lcell_comb \sin_o~16 (
	.dataa(!cordic_y_res_d_16),
	.datab(!cordic_y_res_2c_16),
	.datac(!cordic_x_res_d_16),
	.datad(!cordic_x_res_2c_16),
	.datae(!seg_rot_1),
	.dataf(!seg_rot_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sin_o~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sin_o~16 .extended_lut = "off";
defparam \sin_o~16 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \sin_o~16 .shared_arith = "off";

arriav_lcell_comb \sin_o~17 (
	.dataa(!cordic_y_res_d_17),
	.datab(!cordic_y_res_2c_17),
	.datac(!cordic_x_res_d_17),
	.datad(!cordic_x_res_2c_17),
	.datae(!seg_rot_1),
	.dataf(!seg_rot_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\sin_o~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \sin_o~17 .extended_lut = "off";
defparam \sin_o~17 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \sin_o~17 .shared_arith = "off";

arriav_lcell_comb \cos_o~0 (
	.dataa(!cordic_x_res_d_0),
	.datab(!cordic_x_res_2c_0),
	.datac(!cordic_y_res_2c_0),
	.datad(!cordic_y_res_d_0),
	.datae(!seg_rot_1),
	.dataf(!seg_rot_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cos_o~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cos_o~0 .extended_lut = "off";
defparam \cos_o~0 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \cos_o~0 .shared_arith = "off";

arriav_lcell_comb \cos_o~1 (
	.dataa(!cordic_x_res_d_1),
	.datab(!cordic_x_res_2c_1),
	.datac(!cordic_y_res_2c_1),
	.datad(!cordic_y_res_d_1),
	.datae(!seg_rot_1),
	.dataf(!seg_rot_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cos_o~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cos_o~1 .extended_lut = "off";
defparam \cos_o~1 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \cos_o~1 .shared_arith = "off";

arriav_lcell_comb \cos_o~2 (
	.dataa(!cordic_x_res_d_2),
	.datab(!cordic_x_res_2c_2),
	.datac(!cordic_y_res_2c_2),
	.datad(!cordic_y_res_d_2),
	.datae(!seg_rot_1),
	.dataf(!seg_rot_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cos_o~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cos_o~2 .extended_lut = "off";
defparam \cos_o~2 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \cos_o~2 .shared_arith = "off";

arriav_lcell_comb \cos_o~3 (
	.dataa(!cordic_x_res_d_3),
	.datab(!cordic_x_res_2c_3),
	.datac(!cordic_y_res_2c_3),
	.datad(!cordic_y_res_d_3),
	.datae(!seg_rot_1),
	.dataf(!seg_rot_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cos_o~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cos_o~3 .extended_lut = "off";
defparam \cos_o~3 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \cos_o~3 .shared_arith = "off";

arriav_lcell_comb \cos_o~4 (
	.dataa(!cordic_x_res_d_4),
	.datab(!cordic_x_res_2c_4),
	.datac(!cordic_y_res_2c_4),
	.datad(!cordic_y_res_d_4),
	.datae(!seg_rot_1),
	.dataf(!seg_rot_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cos_o~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cos_o~4 .extended_lut = "off";
defparam \cos_o~4 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \cos_o~4 .shared_arith = "off";

arriav_lcell_comb \cos_o~5 (
	.dataa(!cordic_x_res_d_5),
	.datab(!cordic_x_res_2c_5),
	.datac(!cordic_y_res_2c_5),
	.datad(!cordic_y_res_d_5),
	.datae(!seg_rot_1),
	.dataf(!seg_rot_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cos_o~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cos_o~5 .extended_lut = "off";
defparam \cos_o~5 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \cos_o~5 .shared_arith = "off";

arriav_lcell_comb \cos_o~6 (
	.dataa(!cordic_x_res_d_6),
	.datab(!cordic_x_res_2c_6),
	.datac(!cordic_y_res_2c_6),
	.datad(!cordic_y_res_d_6),
	.datae(!seg_rot_1),
	.dataf(!seg_rot_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cos_o~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cos_o~6 .extended_lut = "off";
defparam \cos_o~6 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \cos_o~6 .shared_arith = "off";

arriav_lcell_comb \cos_o~7 (
	.dataa(!cordic_x_res_d_7),
	.datab(!cordic_x_res_2c_7),
	.datac(!cordic_y_res_2c_7),
	.datad(!cordic_y_res_d_7),
	.datae(!seg_rot_1),
	.dataf(!seg_rot_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cos_o~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cos_o~7 .extended_lut = "off";
defparam \cos_o~7 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \cos_o~7 .shared_arith = "off";

arriav_lcell_comb \cos_o~8 (
	.dataa(!cordic_x_res_d_8),
	.datab(!cordic_x_res_2c_8),
	.datac(!cordic_y_res_2c_8),
	.datad(!cordic_y_res_d_8),
	.datae(!seg_rot_1),
	.dataf(!seg_rot_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cos_o~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cos_o~8 .extended_lut = "off";
defparam \cos_o~8 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \cos_o~8 .shared_arith = "off";

arriav_lcell_comb \cos_o~9 (
	.dataa(!cordic_x_res_d_9),
	.datab(!cordic_x_res_2c_9),
	.datac(!cordic_y_res_2c_9),
	.datad(!cordic_y_res_d_9),
	.datae(!seg_rot_1),
	.dataf(!seg_rot_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cos_o~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cos_o~9 .extended_lut = "off";
defparam \cos_o~9 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \cos_o~9 .shared_arith = "off";

arriav_lcell_comb \cos_o~10 (
	.dataa(!cordic_x_res_d_10),
	.datab(!cordic_x_res_2c_10),
	.datac(!cordic_y_res_2c_10),
	.datad(!cordic_y_res_d_10),
	.datae(!seg_rot_1),
	.dataf(!seg_rot_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cos_o~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cos_o~10 .extended_lut = "off";
defparam \cos_o~10 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \cos_o~10 .shared_arith = "off";

arriav_lcell_comb \cos_o~11 (
	.dataa(!cordic_x_res_d_11),
	.datab(!cordic_x_res_2c_11),
	.datac(!cordic_y_res_2c_11),
	.datad(!cordic_y_res_d_11),
	.datae(!seg_rot_1),
	.dataf(!seg_rot_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cos_o~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cos_o~11 .extended_lut = "off";
defparam \cos_o~11 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \cos_o~11 .shared_arith = "off";

arriav_lcell_comb \cos_o~12 (
	.dataa(!cordic_x_res_d_12),
	.datab(!cordic_x_res_2c_12),
	.datac(!cordic_y_res_2c_12),
	.datad(!cordic_y_res_d_12),
	.datae(!seg_rot_1),
	.dataf(!seg_rot_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cos_o~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cos_o~12 .extended_lut = "off";
defparam \cos_o~12 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \cos_o~12 .shared_arith = "off";

arriav_lcell_comb \cos_o~13 (
	.dataa(!cordic_x_res_d_13),
	.datab(!cordic_x_res_2c_13),
	.datac(!cordic_y_res_2c_13),
	.datad(!cordic_y_res_d_13),
	.datae(!seg_rot_1),
	.dataf(!seg_rot_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cos_o~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cos_o~13 .extended_lut = "off";
defparam \cos_o~13 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \cos_o~13 .shared_arith = "off";

arriav_lcell_comb \cos_o~14 (
	.dataa(!cordic_x_res_d_14),
	.datab(!cordic_x_res_2c_14),
	.datac(!cordic_y_res_2c_14),
	.datad(!cordic_y_res_d_14),
	.datae(!seg_rot_1),
	.dataf(!seg_rot_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cos_o~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cos_o~14 .extended_lut = "off";
defparam \cos_o~14 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \cos_o~14 .shared_arith = "off";

arriav_lcell_comb \cos_o~15 (
	.dataa(!cordic_x_res_d_15),
	.datab(!cordic_x_res_2c_15),
	.datac(!cordic_y_res_2c_15),
	.datad(!cordic_y_res_d_15),
	.datae(!seg_rot_1),
	.dataf(!seg_rot_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cos_o~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cos_o~15 .extended_lut = "off";
defparam \cos_o~15 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \cos_o~15 .shared_arith = "off";

arriav_lcell_comb \cos_o~16 (
	.dataa(!cordic_x_res_d_16),
	.datab(!cordic_x_res_2c_16),
	.datac(!cordic_y_res_2c_16),
	.datad(!cordic_y_res_d_16),
	.datae(!seg_rot_1),
	.dataf(!seg_rot_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cos_o~16_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cos_o~16 .extended_lut = "off";
defparam \cos_o~16 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \cos_o~16 .shared_arith = "off";

arriav_lcell_comb \cos_o~17 (
	.dataa(!cordic_x_res_d_17),
	.datab(!cordic_x_res_2c_17),
	.datac(!cordic_y_res_2c_17),
	.datad(!cordic_y_res_d_17),
	.datae(!seg_rot_1),
	.dataf(!seg_rot_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\cos_o~17_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \cos_o~17 .extended_lut = "off";
defparam \cos_o~17 .lut_mask = 64'h7FFFFFFFFFFF7FFF;
defparam \cos_o~17 .shared_arith = "off";

endmodule

module nco_test_asj_dxx (
	dxxpdo_20,
	dxxpdo_19,
	dxxrv_7,
	dxxrv_6,
	dxxrv_5,
	dxxpdo_18,
	dxxrv_4,
	dxxpdo_17,
	dxxrv_3,
	dxxpdo_16,
	dxxrv_2,
	dxxpdo_15,
	dxxrv_1,
	dxxpdo_14,
	dxxrv_0,
	dxxpdo_13,
	dxxpdo_12,
	dxxpdo_11,
	dxxpdo_10,
	dxxpdo_9,
	dxxpdo_8,
	dxxpdo_7,
	dxxpdo_6,
	dxxpdo_5,
	dxxpdo_4,
	sin_o_0,
	pipeline_dffe_31,
	pipeline_dffe_30,
	pipeline_dffe_29,
	pipeline_dffe_28,
	pipeline_dffe_27,
	pipeline_dffe_26,
	pipeline_dffe_25,
	pipeline_dffe_24,
	pipeline_dffe_23,
	pipeline_dffe_22,
	pipeline_dffe_21,
	pipeline_dffe_20,
	pipeline_dffe_19,
	pipeline_dffe_18,
	pipeline_dffe_17,
	pipeline_dffe_16,
	pipeline_dffe_15,
	pipeline_dffe_14,
	pipeline_dffe_13,
	pipeline_dffe_12,
	pipeline_dffe_11,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	dxxpdo_20;
output 	dxxpdo_19;
input 	dxxrv_7;
input 	dxxrv_6;
input 	dxxrv_5;
output 	dxxpdo_18;
input 	dxxrv_4;
output 	dxxpdo_17;
input 	dxxrv_3;
output 	dxxpdo_16;
input 	dxxrv_2;
output 	dxxpdo_15;
input 	dxxrv_1;
output 	dxxpdo_14;
input 	dxxrv_0;
output 	dxxpdo_13;
output 	dxxpdo_12;
output 	dxxpdo_11;
output 	dxxpdo_10;
output 	dxxpdo_9;
output 	dxxpdo_8;
output 	dxxpdo_7;
output 	dxxpdo_6;
output 	dxxpdo_5;
output 	dxxpdo_4;
input 	sin_o_0;
input 	pipeline_dffe_31;
input 	pipeline_dffe_30;
input 	pipeline_dffe_29;
input 	pipeline_dffe_28;
input 	pipeline_dffe_27;
input 	pipeline_dffe_26;
input 	pipeline_dffe_25;
input 	pipeline_dffe_24;
input 	pipeline_dffe_23;
input 	pipeline_dffe_22;
input 	pipeline_dffe_21;
input 	pipeline_dffe_20;
input 	pipeline_dffe_19;
input 	pipeline_dffe_18;
input 	pipeline_dffe_17;
input 	pipeline_dffe_16;
input 	pipeline_dffe_15;
input 	pipeline_dffe_14;
input 	pipeline_dffe_13;
input 	pipeline_dffe_12;
input 	pipeline_dffe_11;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add0~82_cout ;
wire \Add0~78_cout ;
wire \Add0~74_cout ;
wire \Add0~70_cout ;
wire \Add0~66 ;
wire \Add0~62 ;
wire \Add0~58 ;
wire \Add0~54 ;
wire \Add0~50 ;
wire \Add0~46 ;
wire \Add0~42 ;
wire \Add0~38 ;
wire \Add0~34 ;
wire \Add0~30 ;
wire \Add0~26 ;
wire \Add0~22 ;
wire \Add0~18 ;
wire \Add0~14 ;
wire \Add0~10 ;
wire \Add0~6 ;
wire \Add0~1_sumout ;
wire \phi_dither_out_w[20]~q ;
wire \Add0~5_sumout ;
wire \phi_dither_out_w[19]~q ;
wire \Add0~9_sumout ;
wire \phi_dither_out_w[18]~q ;
wire \Add0~13_sumout ;
wire \phi_dither_out_w[17]~q ;
wire \Add0~17_sumout ;
wire \phi_dither_out_w[16]~q ;
wire \Add0~21_sumout ;
wire \phi_dither_out_w[15]~q ;
wire \Add0~25_sumout ;
wire \phi_dither_out_w[14]~q ;
wire \Add0~29_sumout ;
wire \phi_dither_out_w[13]~q ;
wire \Add0~33_sumout ;
wire \phi_dither_out_w[12]~q ;
wire \Add0~37_sumout ;
wire \phi_dither_out_w[11]~q ;
wire \Add0~41_sumout ;
wire \phi_dither_out_w[10]~q ;
wire \Add0~45_sumout ;
wire \phi_dither_out_w[9]~q ;
wire \Add0~49_sumout ;
wire \phi_dither_out_w[8]~q ;
wire \Add0~53_sumout ;
wire \phi_dither_out_w[7]~q ;
wire \Add0~57_sumout ;
wire \phi_dither_out_w[6]~q ;
wire \Add0~61_sumout ;
wire \phi_dither_out_w[5]~q ;
wire \Add0~65_sumout ;
wire \phi_dither_out_w[4]~q ;


dffeas \dxxpdo[20] (
	.clk(clk),
	.d(\phi_dither_out_w[20]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(dxxpdo_20),
	.prn(vcc));
defparam \dxxpdo[20] .is_wysiwyg = "true";
defparam \dxxpdo[20] .power_up = "low";

dffeas \dxxpdo[19] (
	.clk(clk),
	.d(\phi_dither_out_w[19]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(dxxpdo_19),
	.prn(vcc));
defparam \dxxpdo[19] .is_wysiwyg = "true";
defparam \dxxpdo[19] .power_up = "low";

dffeas \dxxpdo[18] (
	.clk(clk),
	.d(\phi_dither_out_w[18]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(dxxpdo_18),
	.prn(vcc));
defparam \dxxpdo[18] .is_wysiwyg = "true";
defparam \dxxpdo[18] .power_up = "low";

dffeas \dxxpdo[17] (
	.clk(clk),
	.d(\phi_dither_out_w[17]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(dxxpdo_17),
	.prn(vcc));
defparam \dxxpdo[17] .is_wysiwyg = "true";
defparam \dxxpdo[17] .power_up = "low";

dffeas \dxxpdo[16] (
	.clk(clk),
	.d(\phi_dither_out_w[16]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(dxxpdo_16),
	.prn(vcc));
defparam \dxxpdo[16] .is_wysiwyg = "true";
defparam \dxxpdo[16] .power_up = "low";

dffeas \dxxpdo[15] (
	.clk(clk),
	.d(\phi_dither_out_w[15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(dxxpdo_15),
	.prn(vcc));
defparam \dxxpdo[15] .is_wysiwyg = "true";
defparam \dxxpdo[15] .power_up = "low";

dffeas \dxxpdo[14] (
	.clk(clk),
	.d(\phi_dither_out_w[14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(dxxpdo_14),
	.prn(vcc));
defparam \dxxpdo[14] .is_wysiwyg = "true";
defparam \dxxpdo[14] .power_up = "low";

dffeas \dxxpdo[13] (
	.clk(clk),
	.d(\phi_dither_out_w[13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(dxxpdo_13),
	.prn(vcc));
defparam \dxxpdo[13] .is_wysiwyg = "true";
defparam \dxxpdo[13] .power_up = "low";

dffeas \dxxpdo[12] (
	.clk(clk),
	.d(\phi_dither_out_w[12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(dxxpdo_12),
	.prn(vcc));
defparam \dxxpdo[12] .is_wysiwyg = "true";
defparam \dxxpdo[12] .power_up = "low";

dffeas \dxxpdo[11] (
	.clk(clk),
	.d(\phi_dither_out_w[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(dxxpdo_11),
	.prn(vcc));
defparam \dxxpdo[11] .is_wysiwyg = "true";
defparam \dxxpdo[11] .power_up = "low";

dffeas \dxxpdo[10] (
	.clk(clk),
	.d(\phi_dither_out_w[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(dxxpdo_10),
	.prn(vcc));
defparam \dxxpdo[10] .is_wysiwyg = "true";
defparam \dxxpdo[10] .power_up = "low";

dffeas \dxxpdo[9] (
	.clk(clk),
	.d(\phi_dither_out_w[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(dxxpdo_9),
	.prn(vcc));
defparam \dxxpdo[9] .is_wysiwyg = "true";
defparam \dxxpdo[9] .power_up = "low";

dffeas \dxxpdo[8] (
	.clk(clk),
	.d(\phi_dither_out_w[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(dxxpdo_8),
	.prn(vcc));
defparam \dxxpdo[8] .is_wysiwyg = "true";
defparam \dxxpdo[8] .power_up = "low";

dffeas \dxxpdo[7] (
	.clk(clk),
	.d(\phi_dither_out_w[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(dxxpdo_7),
	.prn(vcc));
defparam \dxxpdo[7] .is_wysiwyg = "true";
defparam \dxxpdo[7] .power_up = "low";

dffeas \dxxpdo[6] (
	.clk(clk),
	.d(\phi_dither_out_w[6]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(dxxpdo_6),
	.prn(vcc));
defparam \dxxpdo[6] .is_wysiwyg = "true";
defparam \dxxpdo[6] .power_up = "low";

dffeas \dxxpdo[5] (
	.clk(clk),
	.d(\phi_dither_out_w[5]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(dxxpdo_5),
	.prn(vcc));
defparam \dxxpdo[5] .is_wysiwyg = "true";
defparam \dxxpdo[5] .power_up = "low";

dffeas \dxxpdo[4] (
	.clk(clk),
	.d(\phi_dither_out_w[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(dxxpdo_4),
	.prn(vcc));
defparam \dxxpdo[4] .is_wysiwyg = "true";
defparam \dxxpdo[4] .power_up = "low";

arriav_lcell_comb \Add0~82 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_0),
	.datae(gnd),
	.dataf(!pipeline_dffe_11),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add0~82_cout ),
	.shareout());
defparam \Add0~82 .extended_lut = "off";
defparam \Add0~82 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~82 .shared_arith = "off";

arriav_lcell_comb \Add0~78 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_1),
	.datae(gnd),
	.dataf(!pipeline_dffe_12),
	.datag(gnd),
	.cin(\Add0~82_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add0~78_cout ),
	.shareout());
defparam \Add0~78 .extended_lut = "off";
defparam \Add0~78 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~78 .shared_arith = "off";

arriav_lcell_comb \Add0~74 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_2),
	.datae(gnd),
	.dataf(!pipeline_dffe_13),
	.datag(gnd),
	.cin(\Add0~78_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add0~74_cout ),
	.shareout());
defparam \Add0~74 .extended_lut = "off";
defparam \Add0~74 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~74 .shared_arith = "off";

arriav_lcell_comb \Add0~70 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_3),
	.datae(gnd),
	.dataf(!pipeline_dffe_14),
	.datag(gnd),
	.cin(\Add0~74_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\Add0~70_cout ),
	.shareout());
defparam \Add0~70 .extended_lut = "off";
defparam \Add0~70 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~70 .shared_arith = "off";

arriav_lcell_comb \Add0~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_4),
	.datae(gnd),
	.dataf(!pipeline_dffe_15),
	.datag(gnd),
	.cin(\Add0~70_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~65_sumout ),
	.cout(\Add0~66 ),
	.shareout());
defparam \Add0~65 .extended_lut = "off";
defparam \Add0~65 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~65 .shared_arith = "off";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_5),
	.datae(gnd),
	.dataf(!pipeline_dffe_16),
	.datag(gnd),
	.cin(\Add0~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout());
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~61 .shared_arith = "off";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_6),
	.datae(gnd),
	.dataf(!pipeline_dffe_17),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout());
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~57 .shared_arith = "off";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_7),
	.datae(gnd),
	.dataf(!pipeline_dffe_18),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout());
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~53 .shared_arith = "off";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_7),
	.datae(gnd),
	.dataf(!pipeline_dffe_19),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout());
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~49 .shared_arith = "off";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_7),
	.datae(gnd),
	.dataf(!pipeline_dffe_20),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~45 .shared_arith = "off";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_7),
	.datae(gnd),
	.dataf(!pipeline_dffe_21),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~41 .shared_arith = "off";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_7),
	.datae(gnd),
	.dataf(!pipeline_dffe_22),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~37 .shared_arith = "off";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_7),
	.datae(gnd),
	.dataf(!pipeline_dffe_23),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~33 .shared_arith = "off";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_7),
	.datae(gnd),
	.dataf(!pipeline_dffe_24),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~29 .shared_arith = "off";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_7),
	.datae(gnd),
	.dataf(!pipeline_dffe_25),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~25 .shared_arith = "off";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_7),
	.datae(gnd),
	.dataf(!pipeline_dffe_26),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~21 .shared_arith = "off";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_7),
	.datae(gnd),
	.dataf(!pipeline_dffe_27),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~17 .shared_arith = "off";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_7),
	.datae(gnd),
	.dataf(!pipeline_dffe_28),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~13 .shared_arith = "off";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_7),
	.datae(gnd),
	.dataf(!pipeline_dffe_29),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~9 .shared_arith = "off";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_7),
	.datae(gnd),
	.dataf(!pipeline_dffe_30),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~5 .shared_arith = "off";

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dxxrv_7),
	.datae(gnd),
	.dataf(!pipeline_dffe_31),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~1 .shared_arith = "off";

dffeas \phi_dither_out_w[20] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\phi_dither_out_w[20]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[20] .is_wysiwyg = "true";
defparam \phi_dither_out_w[20] .power_up = "low";

dffeas \phi_dither_out_w[19] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\phi_dither_out_w[19]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[19] .is_wysiwyg = "true";
defparam \phi_dither_out_w[19] .power_up = "low";

dffeas \phi_dither_out_w[18] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\phi_dither_out_w[18]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[18] .is_wysiwyg = "true";
defparam \phi_dither_out_w[18] .power_up = "low";

dffeas \phi_dither_out_w[17] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\phi_dither_out_w[17]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[17] .is_wysiwyg = "true";
defparam \phi_dither_out_w[17] .power_up = "low";

dffeas \phi_dither_out_w[16] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\phi_dither_out_w[16]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[16] .is_wysiwyg = "true";
defparam \phi_dither_out_w[16] .power_up = "low";

dffeas \phi_dither_out_w[15] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\phi_dither_out_w[15]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[15] .is_wysiwyg = "true";
defparam \phi_dither_out_w[15] .power_up = "low";

dffeas \phi_dither_out_w[14] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\phi_dither_out_w[14]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[14] .is_wysiwyg = "true";
defparam \phi_dither_out_w[14] .power_up = "low";

dffeas \phi_dither_out_w[13] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\phi_dither_out_w[13]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[13] .is_wysiwyg = "true";
defparam \phi_dither_out_w[13] .power_up = "low";

dffeas \phi_dither_out_w[12] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\phi_dither_out_w[12]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[12] .is_wysiwyg = "true";
defparam \phi_dither_out_w[12] .power_up = "low";

dffeas \phi_dither_out_w[11] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\phi_dither_out_w[11]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[11] .is_wysiwyg = "true";
defparam \phi_dither_out_w[11] .power_up = "low";

dffeas \phi_dither_out_w[10] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\phi_dither_out_w[10]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[10] .is_wysiwyg = "true";
defparam \phi_dither_out_w[10] .power_up = "low";

dffeas \phi_dither_out_w[9] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\phi_dither_out_w[9]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[9] .is_wysiwyg = "true";
defparam \phi_dither_out_w[9] .power_up = "low";

dffeas \phi_dither_out_w[8] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\phi_dither_out_w[8]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[8] .is_wysiwyg = "true";
defparam \phi_dither_out_w[8] .power_up = "low";

dffeas \phi_dither_out_w[7] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\phi_dither_out_w[7]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[7] .is_wysiwyg = "true";
defparam \phi_dither_out_w[7] .power_up = "low";

dffeas \phi_dither_out_w[6] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\phi_dither_out_w[6]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[6] .is_wysiwyg = "true";
defparam \phi_dither_out_w[6] .power_up = "low";

dffeas \phi_dither_out_w[5] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\phi_dither_out_w[5]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[5] .is_wysiwyg = "true";
defparam \phi_dither_out_w[5] .power_up = "low";

dffeas \phi_dither_out_w[4] (
	.clk(clk),
	.d(\Add0~65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\phi_dither_out_w[4]~q ),
	.prn(vcc));
defparam \phi_dither_out_w[4] .is_wysiwyg = "true";
defparam \phi_dither_out_w[4] .power_up = "low";

endmodule

module nco_test_asj_dxx_g (
	dxxrv_7,
	dxxrv_6,
	dxxrv_5,
	dxxrv_4,
	dxxrv_3,
	dxxrv_2,
	dxxrv_1,
	dxxrv_0,
	sin_o_0,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	dxxrv_7;
output 	dxxrv_6;
output 	dxxrv_5;
output 	dxxrv_4;
output 	dxxrv_3;
output 	dxxrv_2;
output 	dxxrv_1;
output 	dxxrv_0;
input 	sin_o_0;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \lsfr_reg~9_combout ;
wire \lsfr_reg[0]~q ;
wire \lsfr_reg[1]~q ;
wire \lsfr_reg~8_combout ;
wire \lsfr_reg[2]~q ;
wire \lsfr_reg~7_combout ;
wire \lsfr_reg[3]~q ;
wire \lsfr_reg~6_combout ;
wire \lsfr_reg[4]~q ;
wire \lsfr_reg[5]~q ;
wire \lsfr_reg~5_combout ;
wire \lsfr_reg[6]~q ;
wire \lsfr_reg~4_combout ;
wire \lsfr_reg[7]~q ;
wire \lsfr_reg[8]~q ;
wire \lsfr_reg~3_combout ;
wire \lsfr_reg[9]~q ;
wire \lsfr_reg[10]~q ;
wire \lsfr_reg~2_combout ;
wire \lsfr_reg[11]~q ;
wire \lsfr_reg~1_combout ;
wire \lsfr_reg[12]~q ;
wire \lsfr_reg[13]~q ;
wire \lsfr_reg[14]~q ;
wire \lsfr_reg~0_combout ;
wire \lsfr_reg[15]~q ;
wire \Add0~30 ;
wire \Add0~26 ;
wire \Add0~22 ;
wire \Add0~18 ;
wire \Add0~14 ;
wire \Add0~10 ;
wire \Add0~6 ;
wire \Add0~1_sumout ;
wire \Add0~5_sumout ;
wire \Add0~9_sumout ;
wire \Add0~13_sumout ;
wire \Add0~17_sumout ;
wire \Add0~21_sumout ;
wire \Add0~25_sumout ;
wire \Add0~29_sumout ;


dffeas \dxxrv[7] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(dxxrv_7),
	.prn(vcc));
defparam \dxxrv[7] .is_wysiwyg = "true";
defparam \dxxrv[7] .power_up = "low";

dffeas \dxxrv[6] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(dxxrv_6),
	.prn(vcc));
defparam \dxxrv[6] .is_wysiwyg = "true";
defparam \dxxrv[6] .power_up = "low";

dffeas \dxxrv[5] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(dxxrv_5),
	.prn(vcc));
defparam \dxxrv[5] .is_wysiwyg = "true";
defparam \dxxrv[5] .power_up = "low";

dffeas \dxxrv[4] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(dxxrv_4),
	.prn(vcc));
defparam \dxxrv[4] .is_wysiwyg = "true";
defparam \dxxrv[4] .power_up = "low";

dffeas \dxxrv[3] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(dxxrv_3),
	.prn(vcc));
defparam \dxxrv[3] .is_wysiwyg = "true";
defparam \dxxrv[3] .power_up = "low";

dffeas \dxxrv[2] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(dxxrv_2),
	.prn(vcc));
defparam \dxxrv[2] .is_wysiwyg = "true";
defparam \dxxrv[2] .power_up = "low";

dffeas \dxxrv[1] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(dxxrv_1),
	.prn(vcc));
defparam \dxxrv[1] .is_wysiwyg = "true";
defparam \dxxrv[1] .power_up = "low";

dffeas \dxxrv[0] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(dxxrv_0),
	.prn(vcc));
defparam \dxxrv[0] .is_wysiwyg = "true";
defparam \dxxrv[0] .power_up = "low";

arriav_lcell_comb \lsfr_reg~9 (
	.dataa(!\lsfr_reg[15]~q ),
	.datab(!\lsfr_reg[14]~q ),
	.datac(!\lsfr_reg[12]~q ),
	.datad(!\lsfr_reg[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg~9 .extended_lut = "off";
defparam \lsfr_reg~9 .lut_mask = 64'h6996699669966996;
defparam \lsfr_reg~9 .shared_arith = "off";

dffeas \lsfr_reg[0] (
	.clk(clk),
	.d(\lsfr_reg~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(!reset_n),
	.ena(sin_o_0),
	.q(\lsfr_reg[0]~q ),
	.prn(vcc));
defparam \lsfr_reg[0] .is_wysiwyg = "true";
defparam \lsfr_reg[0] .power_up = "low";

dffeas \lsfr_reg[1] (
	.clk(clk),
	.d(\lsfr_reg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\lsfr_reg[1]~q ),
	.prn(vcc));
defparam \lsfr_reg[1] .is_wysiwyg = "true";
defparam \lsfr_reg[1] .power_up = "low";

arriav_lcell_comb \lsfr_reg~8 (
	.dataa(!reset_n),
	.datab(!\lsfr_reg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg~8 .extended_lut = "off";
defparam \lsfr_reg~8 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \lsfr_reg~8 .shared_arith = "off";

dffeas \lsfr_reg[2] (
	.clk(clk),
	.d(\lsfr_reg~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\lsfr_reg[2]~q ),
	.prn(vcc));
defparam \lsfr_reg[2] .is_wysiwyg = "true";
defparam \lsfr_reg[2] .power_up = "low";

arriav_lcell_comb \lsfr_reg~7 (
	.dataa(!reset_n),
	.datab(!\lsfr_reg[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg~7 .extended_lut = "off";
defparam \lsfr_reg~7 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \lsfr_reg~7 .shared_arith = "off";

dffeas \lsfr_reg[3] (
	.clk(clk),
	.d(\lsfr_reg~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\lsfr_reg[3]~q ),
	.prn(vcc));
defparam \lsfr_reg[3] .is_wysiwyg = "true";
defparam \lsfr_reg[3] .power_up = "low";

arriav_lcell_comb \lsfr_reg~6 (
	.dataa(!reset_n),
	.datab(!\lsfr_reg[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg~6 .extended_lut = "off";
defparam \lsfr_reg~6 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \lsfr_reg~6 .shared_arith = "off";

dffeas \lsfr_reg[4] (
	.clk(clk),
	.d(\lsfr_reg~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\lsfr_reg[4]~q ),
	.prn(vcc));
defparam \lsfr_reg[4] .is_wysiwyg = "true";
defparam \lsfr_reg[4] .power_up = "low";

dffeas \lsfr_reg[5] (
	.clk(clk),
	.d(\lsfr_reg[4]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\lsfr_reg[5]~q ),
	.prn(vcc));
defparam \lsfr_reg[5] .is_wysiwyg = "true";
defparam \lsfr_reg[5] .power_up = "low";

arriav_lcell_comb \lsfr_reg~5 (
	.dataa(!reset_n),
	.datab(!\lsfr_reg[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg~5 .extended_lut = "off";
defparam \lsfr_reg~5 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \lsfr_reg~5 .shared_arith = "off";

dffeas \lsfr_reg[6] (
	.clk(clk),
	.d(\lsfr_reg~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\lsfr_reg[6]~q ),
	.prn(vcc));
defparam \lsfr_reg[6] .is_wysiwyg = "true";
defparam \lsfr_reg[6] .power_up = "low";

arriav_lcell_comb \lsfr_reg~4 (
	.dataa(!reset_n),
	.datab(!\lsfr_reg[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg~4 .extended_lut = "off";
defparam \lsfr_reg~4 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \lsfr_reg~4 .shared_arith = "off";

dffeas \lsfr_reg[7] (
	.clk(clk),
	.d(\lsfr_reg~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\lsfr_reg[7]~q ),
	.prn(vcc));
defparam \lsfr_reg[7] .is_wysiwyg = "true";
defparam \lsfr_reg[7] .power_up = "low";

dffeas \lsfr_reg[8] (
	.clk(clk),
	.d(\lsfr_reg[7]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\lsfr_reg[8]~q ),
	.prn(vcc));
defparam \lsfr_reg[8] .is_wysiwyg = "true";
defparam \lsfr_reg[8] .power_up = "low";

arriav_lcell_comb \lsfr_reg~3 (
	.dataa(!reset_n),
	.datab(!\lsfr_reg[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg~3 .extended_lut = "off";
defparam \lsfr_reg~3 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \lsfr_reg~3 .shared_arith = "off";

dffeas \lsfr_reg[9] (
	.clk(clk),
	.d(\lsfr_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\lsfr_reg[9]~q ),
	.prn(vcc));
defparam \lsfr_reg[9] .is_wysiwyg = "true";
defparam \lsfr_reg[9] .power_up = "low";

dffeas \lsfr_reg[10] (
	.clk(clk),
	.d(\lsfr_reg[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\lsfr_reg[10]~q ),
	.prn(vcc));
defparam \lsfr_reg[10] .is_wysiwyg = "true";
defparam \lsfr_reg[10] .power_up = "low";

arriav_lcell_comb \lsfr_reg~2 (
	.dataa(!reset_n),
	.datab(!\lsfr_reg[10]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg~2 .extended_lut = "off";
defparam \lsfr_reg~2 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \lsfr_reg~2 .shared_arith = "off";

dffeas \lsfr_reg[11] (
	.clk(clk),
	.d(\lsfr_reg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\lsfr_reg[11]~q ),
	.prn(vcc));
defparam \lsfr_reg[11] .is_wysiwyg = "true";
defparam \lsfr_reg[11] .power_up = "low";

arriav_lcell_comb \lsfr_reg~1 (
	.dataa(!reset_n),
	.datab(!\lsfr_reg[11]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg~1 .extended_lut = "off";
defparam \lsfr_reg~1 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \lsfr_reg~1 .shared_arith = "off";

dffeas \lsfr_reg[12] (
	.clk(clk),
	.d(\lsfr_reg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\lsfr_reg[12]~q ),
	.prn(vcc));
defparam \lsfr_reg[12] .is_wysiwyg = "true";
defparam \lsfr_reg[12] .power_up = "low";

dffeas \lsfr_reg[13] (
	.clk(clk),
	.d(\lsfr_reg[12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\lsfr_reg[13]~q ),
	.prn(vcc));
defparam \lsfr_reg[13] .is_wysiwyg = "true";
defparam \lsfr_reg[13] .power_up = "low";

dffeas \lsfr_reg[14] (
	.clk(clk),
	.d(\lsfr_reg[13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\lsfr_reg[14]~q ),
	.prn(vcc));
defparam \lsfr_reg[14] .is_wysiwyg = "true";
defparam \lsfr_reg[14] .power_up = "low";

arriav_lcell_comb \lsfr_reg~0 (
	.dataa(!reset_n),
	.datab(!\lsfr_reg[14]~q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\lsfr_reg~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \lsfr_reg~0 .extended_lut = "off";
defparam \lsfr_reg~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \lsfr_reg~0 .shared_arith = "off";

dffeas \lsfr_reg[15] (
	.clk(clk),
	.d(\lsfr_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\lsfr_reg[15]~q ),
	.prn(vcc));
defparam \lsfr_reg[15] .is_wysiwyg = "true";
defparam \lsfr_reg[15] .power_up = "low";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\lsfr_reg[8]~q ),
	.datae(gnd),
	.dataf(!\lsfr_reg[15]~q ),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~29 .shared_arith = "off";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\lsfr_reg[9]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h00000000000000FF;
defparam \Add0~25 .shared_arith = "off";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\lsfr_reg[10]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h00000000000000FF;
defparam \Add0~21 .shared_arith = "off";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\lsfr_reg[11]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h00000000000000FF;
defparam \Add0~17 .shared_arith = "off";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\lsfr_reg[12]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h00000000000000FF;
defparam \Add0~13 .shared_arith = "off";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\lsfr_reg[13]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h00000000000000FF;
defparam \Add0~9 .shared_arith = "off";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\lsfr_reg[14]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h00000000000000FF;
defparam \Add0~5 .shared_arith = "off";

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!\lsfr_reg[15]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h00000000000000FF;
defparam \Add0~1 .shared_arith = "off";

endmodule

module nco_test_asj_nco_isdr (
	data_ready1,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	data_ready1;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \lpm_counter_component|auto_generated|counter_reg_bit[2]~q ;
wire \lpm_counter_component|auto_generated|counter_reg_bit[1]~q ;
wire \lpm_counter_component|auto_generated|counter_reg_bit[0]~q ;
wire \lpm_counter_component|auto_generated|counter_reg_bit[5]~q ;
wire \lpm_counter_component|auto_generated|counter_reg_bit[4]~q ;
wire \lpm_counter_component|auto_generated|counter_reg_bit[3]~q ;
wire \always0~0_combout ;
wire \data_ready~0_combout ;


nco_test_lpm_counter_1 lpm_counter_component(
	.counter_reg_bit_2(\lpm_counter_component|auto_generated|counter_reg_bit[2]~q ),
	.counter_reg_bit_1(\lpm_counter_component|auto_generated|counter_reg_bit[1]~q ),
	.counter_reg_bit_0(\lpm_counter_component|auto_generated|counter_reg_bit[0]~q ),
	.counter_reg_bit_5(\lpm_counter_component|auto_generated|counter_reg_bit[5]~q ),
	.counter_reg_bit_4(\lpm_counter_component|auto_generated|counter_reg_bit[4]~q ),
	.counter_reg_bit_3(\lpm_counter_component|auto_generated|counter_reg_bit[3]~q ),
	.clock(clk),
	.sclr(reset_n),
	.clken(clken));

dffeas data_ready(
	.clk(clk),
	.d(\data_ready~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(vcc),
	.q(data_ready1),
	.prn(vcc));
defparam data_ready.is_wysiwyg = "true";
defparam data_ready.power_up = "low";

arriav_lcell_comb \always0~0 (
	.dataa(!clken),
	.datab(!\lpm_counter_component|auto_generated|counter_reg_bit[5]~q ),
	.datac(!\lpm_counter_component|auto_generated|counter_reg_bit[4]~q ),
	.datad(!\lpm_counter_component|auto_generated|counter_reg_bit[3]~q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\always0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \always0~0 .extended_lut = "off";
defparam \always0~0 .lut_mask = 64'hF7FFF7FFF7FFF7FF;
defparam \always0~0 .shared_arith = "off";

arriav_lcell_comb \data_ready~0 (
	.dataa(!data_ready1),
	.datab(!\lpm_counter_component|auto_generated|counter_reg_bit[2]~q ),
	.datac(!\lpm_counter_component|auto_generated|counter_reg_bit[1]~q ),
	.datad(!\lpm_counter_component|auto_generated|counter_reg_bit[0]~q ),
	.datae(!\always0~0_combout ),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\data_ready~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \data_ready~0 .extended_lut = "off";
defparam \data_ready~0 .lut_mask = 64'hFFDFFFFFFFDFFFFF;
defparam \data_ready~0 .shared_arith = "off";

endmodule

module nco_test_lpm_counter_1 (
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	clock,
	sclr,
	clken)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
input 	clock;
input 	sclr;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_cntr_0ei auto_generated(
	.counter_reg_bit_2(counter_reg_bit_2),
	.counter_reg_bit_1(counter_reg_bit_1),
	.counter_reg_bit_0(counter_reg_bit_0),
	.counter_reg_bit_5(counter_reg_bit_5),
	.counter_reg_bit_4(counter_reg_bit_4),
	.counter_reg_bit_3(counter_reg_bit_3),
	.clock(clock),
	.sclr(sclr),
	.clken(clken));

endmodule

module nco_test_cntr_0ei (
	counter_reg_bit_2,
	counter_reg_bit_1,
	counter_reg_bit_0,
	counter_reg_bit_5,
	counter_reg_bit_4,
	counter_reg_bit_3,
	clock,
	sclr,
	clken)/* synthesis synthesis_greybox=1 */;
output 	counter_reg_bit_2;
output 	counter_reg_bit_1;
output 	counter_reg_bit_0;
output 	counter_reg_bit_5;
output 	counter_reg_bit_4;
output 	counter_reg_bit_3;
input 	clock;
input 	sclr;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \counter_comb_bita0~COUT ;
wire \counter_comb_bita1~COUT ;
wire \counter_comb_bita2~sumout ;
wire \counter_comb_bita1~sumout ;
wire \counter_comb_bita0~sumout ;
wire \counter_comb_bita2~COUT ;
wire \counter_comb_bita3~COUT ;
wire \counter_comb_bita4~COUT ;
wire \counter_comb_bita5~sumout ;
wire \counter_comb_bita4~sumout ;
wire \counter_comb_bita3~sumout ;


dffeas \counter_reg_bit[2] (
	.clk(clock),
	.d(\counter_comb_bita2~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sclr),
	.sload(gnd),
	.ena(clken),
	.q(counter_reg_bit_2),
	.prn(vcc));
defparam \counter_reg_bit[2] .is_wysiwyg = "true";
defparam \counter_reg_bit[2] .power_up = "low";

dffeas \counter_reg_bit[1] (
	.clk(clock),
	.d(\counter_comb_bita1~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sclr),
	.sload(gnd),
	.ena(clken),
	.q(counter_reg_bit_1),
	.prn(vcc));
defparam \counter_reg_bit[1] .is_wysiwyg = "true";
defparam \counter_reg_bit[1] .power_up = "low";

dffeas \counter_reg_bit[0] (
	.clk(clock),
	.d(\counter_comb_bita0~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sclr),
	.sload(gnd),
	.ena(clken),
	.q(counter_reg_bit_0),
	.prn(vcc));
defparam \counter_reg_bit[0] .is_wysiwyg = "true";
defparam \counter_reg_bit[0] .power_up = "low";

dffeas \counter_reg_bit[5] (
	.clk(clock),
	.d(\counter_comb_bita5~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sclr),
	.sload(gnd),
	.ena(clken),
	.q(counter_reg_bit_5),
	.prn(vcc));
defparam \counter_reg_bit[5] .is_wysiwyg = "true";
defparam \counter_reg_bit[5] .power_up = "low";

dffeas \counter_reg_bit[4] (
	.clk(clock),
	.d(\counter_comb_bita4~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sclr),
	.sload(gnd),
	.ena(clken),
	.q(counter_reg_bit_4),
	.prn(vcc));
defparam \counter_reg_bit[4] .is_wysiwyg = "true";
defparam \counter_reg_bit[4] .power_up = "low";

dffeas \counter_reg_bit[3] (
	.clk(clock),
	.d(\counter_comb_bita3~sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!sclr),
	.sload(gnd),
	.ena(clken),
	.q(counter_reg_bit_3),
	.prn(vcc));
defparam \counter_reg_bit[3] .is_wysiwyg = "true";
defparam \counter_reg_bit[3] .power_up = "low";

arriav_lcell_comb counter_comb_bita0(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita0~sumout ),
	.cout(\counter_comb_bita0~COUT ),
	.shareout());
defparam counter_comb_bita0.extended_lut = "off";
defparam counter_comb_bita0.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita0.shared_arith = "off";

arriav_lcell_comb counter_comb_bita1(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita0~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita1~sumout ),
	.cout(\counter_comb_bita1~COUT ),
	.shareout());
defparam counter_comb_bita1.extended_lut = "off";
defparam counter_comb_bita1.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita1.shared_arith = "off";

arriav_lcell_comb counter_comb_bita2(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita1~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita2~sumout ),
	.cout(\counter_comb_bita2~COUT ),
	.shareout());
defparam counter_comb_bita2.extended_lut = "off";
defparam counter_comb_bita2.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita2.shared_arith = "off";

arriav_lcell_comb counter_comb_bita3(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita2~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita3~sumout ),
	.cout(\counter_comb_bita3~COUT ),
	.shareout());
defparam counter_comb_bita3.extended_lut = "off";
defparam counter_comb_bita3.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita3.shared_arith = "off";

arriav_lcell_comb counter_comb_bita4(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita3~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita4~sumout ),
	.cout(\counter_comb_bita4~COUT ),
	.shareout());
defparam counter_comb_bita4.extended_lut = "off";
defparam counter_comb_bita4.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita4.shared_arith = "off";

arriav_lcell_comb counter_comb_bita5(
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!counter_reg_bit_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\counter_comb_bita4~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\counter_comb_bita5~sumout ),
	.cout(),
	.shareout());
defparam counter_comb_bita5.extended_lut = "off";
defparam counter_comb_bita5.lut_mask = 64'h00000000000000FF;
defparam counter_comb_bita5.shared_arith = "off";

endmodule

module nco_test_cord_2c (
	cordic_y_res_d_0,
	cordic_y_res_2c_0,
	cordic_x_res_d_0,
	cordic_x_res_2c_0,
	cordic_y_res_d_1,
	cordic_y_res_2c_1,
	cordic_x_res_d_1,
	cordic_x_res_2c_1,
	cordic_y_res_d_2,
	cordic_y_res_2c_2,
	cordic_x_res_d_2,
	cordic_x_res_2c_2,
	cordic_y_res_d_3,
	cordic_y_res_2c_3,
	cordic_x_res_d_3,
	cordic_x_res_2c_3,
	cordic_y_res_d_4,
	cordic_y_res_2c_4,
	cordic_x_res_d_4,
	cordic_x_res_2c_4,
	cordic_y_res_d_5,
	cordic_y_res_2c_5,
	cordic_x_res_d_5,
	cordic_x_res_2c_5,
	cordic_y_res_d_6,
	cordic_y_res_2c_6,
	cordic_x_res_d_6,
	cordic_x_res_2c_6,
	cordic_y_res_d_7,
	cordic_y_res_2c_7,
	cordic_x_res_d_7,
	cordic_x_res_2c_7,
	cordic_y_res_d_8,
	cordic_y_res_2c_8,
	cordic_x_res_d_8,
	cordic_x_res_2c_8,
	cordic_y_res_d_9,
	cordic_y_res_2c_9,
	cordic_x_res_d_9,
	cordic_x_res_2c_9,
	cordic_y_res_d_10,
	cordic_y_res_2c_10,
	cordic_x_res_d_10,
	cordic_x_res_2c_10,
	cordic_y_res_d_11,
	cordic_y_res_2c_11,
	cordic_x_res_d_11,
	cordic_x_res_2c_11,
	cordic_y_res_d_12,
	cordic_y_res_2c_12,
	cordic_x_res_d_12,
	cordic_x_res_2c_12,
	cordic_y_res_d_13,
	cordic_y_res_2c_13,
	cordic_x_res_d_13,
	cordic_x_res_2c_13,
	cordic_y_res_d_14,
	cordic_y_res_2c_14,
	cordic_x_res_d_14,
	cordic_x_res_2c_14,
	cordic_y_res_d_15,
	cordic_y_res_2c_15,
	cordic_x_res_d_15,
	cordic_x_res_2c_15,
	cordic_y_res_d_16,
	cordic_y_res_2c_16,
	cordic_x_res_d_16,
	cordic_x_res_2c_16,
	cordic_y_res_d_17,
	cordic_y_res_2c_17,
	cordic_x_res_d_17,
	cordic_x_res_2c_17,
	sin_o_0,
	pipeline_dffe_0,
	dffe1,
	pipeline_dffe_1,
	dffe2,
	pipeline_dffe_2,
	dffe3,
	pipeline_dffe_3,
	dffe4,
	pipeline_dffe_4,
	dffe5,
	pipeline_dffe_5,
	dffe6,
	pipeline_dffe_6,
	dffe7,
	pipeline_dffe_7,
	dffe8,
	pipeline_dffe_8,
	dffe9,
	pipeline_dffe_9,
	dffe10,
	pipeline_dffe_10,
	dffe11,
	pipeline_dffe_11,
	dffe12,
	pipeline_dffe_12,
	dffe13,
	pipeline_dffe_13,
	dffe14,
	pipeline_dffe_14,
	dffe15,
	pipeline_dffe_15,
	dffe16,
	pipeline_dffe_16,
	dffe17,
	pipeline_dffe_17,
	dffe18,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	cordic_y_res_d_0;
output 	cordic_y_res_2c_0;
output 	cordic_x_res_d_0;
output 	cordic_x_res_2c_0;
output 	cordic_y_res_d_1;
output 	cordic_y_res_2c_1;
output 	cordic_x_res_d_1;
output 	cordic_x_res_2c_1;
output 	cordic_y_res_d_2;
output 	cordic_y_res_2c_2;
output 	cordic_x_res_d_2;
output 	cordic_x_res_2c_2;
output 	cordic_y_res_d_3;
output 	cordic_y_res_2c_3;
output 	cordic_x_res_d_3;
output 	cordic_x_res_2c_3;
output 	cordic_y_res_d_4;
output 	cordic_y_res_2c_4;
output 	cordic_x_res_d_4;
output 	cordic_x_res_2c_4;
output 	cordic_y_res_d_5;
output 	cordic_y_res_2c_5;
output 	cordic_x_res_d_5;
output 	cordic_x_res_2c_5;
output 	cordic_y_res_d_6;
output 	cordic_y_res_2c_6;
output 	cordic_x_res_d_6;
output 	cordic_x_res_2c_6;
output 	cordic_y_res_d_7;
output 	cordic_y_res_2c_7;
output 	cordic_x_res_d_7;
output 	cordic_x_res_2c_7;
output 	cordic_y_res_d_8;
output 	cordic_y_res_2c_8;
output 	cordic_x_res_d_8;
output 	cordic_x_res_2c_8;
output 	cordic_y_res_d_9;
output 	cordic_y_res_2c_9;
output 	cordic_x_res_d_9;
output 	cordic_x_res_2c_9;
output 	cordic_y_res_d_10;
output 	cordic_y_res_2c_10;
output 	cordic_x_res_d_10;
output 	cordic_x_res_2c_10;
output 	cordic_y_res_d_11;
output 	cordic_y_res_2c_11;
output 	cordic_x_res_d_11;
output 	cordic_x_res_2c_11;
output 	cordic_y_res_d_12;
output 	cordic_y_res_2c_12;
output 	cordic_x_res_d_12;
output 	cordic_x_res_2c_12;
output 	cordic_y_res_d_13;
output 	cordic_y_res_2c_13;
output 	cordic_x_res_d_13;
output 	cordic_x_res_2c_13;
output 	cordic_y_res_d_14;
output 	cordic_y_res_2c_14;
output 	cordic_x_res_d_14;
output 	cordic_x_res_2c_14;
output 	cordic_y_res_d_15;
output 	cordic_y_res_2c_15;
output 	cordic_x_res_d_15;
output 	cordic_x_res_2c_15;
output 	cordic_y_res_d_16;
output 	cordic_y_res_2c_16;
output 	cordic_x_res_d_16;
output 	cordic_x_res_2c_16;
output 	cordic_y_res_d_17;
output 	cordic_y_res_2c_17;
output 	cordic_x_res_d_17;
output 	cordic_x_res_2c_17;
input 	sin_o_0;
input 	pipeline_dffe_0;
input 	dffe1;
input 	pipeline_dffe_1;
input 	dffe2;
input 	pipeline_dffe_2;
input 	dffe3;
input 	pipeline_dffe_3;
input 	dffe4;
input 	pipeline_dffe_4;
input 	dffe5;
input 	pipeline_dffe_5;
input 	dffe6;
input 	pipeline_dffe_6;
input 	dffe7;
input 	pipeline_dffe_7;
input 	dffe8;
input 	pipeline_dffe_8;
input 	dffe9;
input 	pipeline_dffe_9;
input 	dffe10;
input 	pipeline_dffe_10;
input 	dffe11;
input 	pipeline_dffe_11;
input 	dffe12;
input 	pipeline_dffe_12;
input 	dffe13;
input 	pipeline_dffe_13;
input 	dffe14;
input 	pipeline_dffe_14;
input 	dffe15;
input 	pipeline_dffe_15;
input 	dffe16;
input 	pipeline_dffe_16;
input 	dffe17;
input 	pipeline_dffe_17;
input 	dffe18;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Add1~1_sumout ;
wire \Add0~1_sumout ;
wire \Add1~2 ;
wire \Add1~5_sumout ;
wire \Add0~2 ;
wire \Add0~5_sumout ;
wire \Add1~6 ;
wire \Add1~9_sumout ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \Add1~10 ;
wire \Add1~13_sumout ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \Add1~14 ;
wire \Add1~17_sumout ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \Add1~18 ;
wire \Add1~21_sumout ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \Add1~22 ;
wire \Add1~25_sumout ;
wire \Add0~22 ;
wire \Add0~25_sumout ;
wire \Add1~26 ;
wire \Add1~29_sumout ;
wire \Add0~26 ;
wire \Add0~29_sumout ;
wire \Add1~30 ;
wire \Add1~33_sumout ;
wire \Add0~30 ;
wire \Add0~33_sumout ;
wire \Add1~34 ;
wire \Add1~37_sumout ;
wire \Add0~34 ;
wire \Add0~37_sumout ;
wire \Add1~38 ;
wire \Add1~41_sumout ;
wire \Add0~38 ;
wire \Add0~41_sumout ;
wire \Add1~42 ;
wire \Add1~45_sumout ;
wire \Add0~42 ;
wire \Add0~45_sumout ;
wire \Add1~46 ;
wire \Add1~49_sumout ;
wire \Add0~46 ;
wire \Add0~49_sumout ;
wire \Add1~50 ;
wire \Add1~53_sumout ;
wire \Add0~50 ;
wire \Add0~53_sumout ;
wire \Add1~54 ;
wire \Add1~57_sumout ;
wire \Add0~54 ;
wire \Add0~57_sumout ;
wire \Add1~58 ;
wire \Add1~61_sumout ;
wire \Add0~58 ;
wire \Add0~61_sumout ;
wire \Add1~62 ;
wire \Add1~65_sumout ;
wire \Add0~62 ;
wire \Add0~65_sumout ;
wire \Add1~66 ;
wire \Add1~69_sumout ;
wire \Add0~66 ;
wire \Add0~69_sumout ;


dffeas \cordic_y_res_d[0] (
	.clk(clk),
	.d(pipeline_dffe_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_y_res_d_0),
	.prn(vcc));
defparam \cordic_y_res_d[0] .is_wysiwyg = "true";
defparam \cordic_y_res_d[0] .power_up = "low";

dffeas \cordic_y_res_2c[0] (
	.clk(clk),
	.d(\Add1~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_y_res_2c_0),
	.prn(vcc));
defparam \cordic_y_res_2c[0] .is_wysiwyg = "true";
defparam \cordic_y_res_2c[0] .power_up = "low";

dffeas \cordic_x_res_d[0] (
	.clk(clk),
	.d(dffe1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_x_res_d_0),
	.prn(vcc));
defparam \cordic_x_res_d[0] .is_wysiwyg = "true";
defparam \cordic_x_res_d[0] .power_up = "low";

dffeas \cordic_x_res_2c[0] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_x_res_2c_0),
	.prn(vcc));
defparam \cordic_x_res_2c[0] .is_wysiwyg = "true";
defparam \cordic_x_res_2c[0] .power_up = "low";

dffeas \cordic_y_res_d[1] (
	.clk(clk),
	.d(pipeline_dffe_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_y_res_d_1),
	.prn(vcc));
defparam \cordic_y_res_d[1] .is_wysiwyg = "true";
defparam \cordic_y_res_d[1] .power_up = "low";

dffeas \cordic_y_res_2c[1] (
	.clk(clk),
	.d(\Add1~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_y_res_2c_1),
	.prn(vcc));
defparam \cordic_y_res_2c[1] .is_wysiwyg = "true";
defparam \cordic_y_res_2c[1] .power_up = "low";

dffeas \cordic_x_res_d[1] (
	.clk(clk),
	.d(dffe2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_x_res_d_1),
	.prn(vcc));
defparam \cordic_x_res_d[1] .is_wysiwyg = "true";
defparam \cordic_x_res_d[1] .power_up = "low";

dffeas \cordic_x_res_2c[1] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_x_res_2c_1),
	.prn(vcc));
defparam \cordic_x_res_2c[1] .is_wysiwyg = "true";
defparam \cordic_x_res_2c[1] .power_up = "low";

dffeas \cordic_y_res_d[2] (
	.clk(clk),
	.d(pipeline_dffe_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_y_res_d_2),
	.prn(vcc));
defparam \cordic_y_res_d[2] .is_wysiwyg = "true";
defparam \cordic_y_res_d[2] .power_up = "low";

dffeas \cordic_y_res_2c[2] (
	.clk(clk),
	.d(\Add1~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_y_res_2c_2),
	.prn(vcc));
defparam \cordic_y_res_2c[2] .is_wysiwyg = "true";
defparam \cordic_y_res_2c[2] .power_up = "low";

dffeas \cordic_x_res_d[2] (
	.clk(clk),
	.d(dffe3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_x_res_d_2),
	.prn(vcc));
defparam \cordic_x_res_d[2] .is_wysiwyg = "true";
defparam \cordic_x_res_d[2] .power_up = "low";

dffeas \cordic_x_res_2c[2] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_x_res_2c_2),
	.prn(vcc));
defparam \cordic_x_res_2c[2] .is_wysiwyg = "true";
defparam \cordic_x_res_2c[2] .power_up = "low";

dffeas \cordic_y_res_d[3] (
	.clk(clk),
	.d(pipeline_dffe_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_y_res_d_3),
	.prn(vcc));
defparam \cordic_y_res_d[3] .is_wysiwyg = "true";
defparam \cordic_y_res_d[3] .power_up = "low";

dffeas \cordic_y_res_2c[3] (
	.clk(clk),
	.d(\Add1~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_y_res_2c_3),
	.prn(vcc));
defparam \cordic_y_res_2c[3] .is_wysiwyg = "true";
defparam \cordic_y_res_2c[3] .power_up = "low";

dffeas \cordic_x_res_d[3] (
	.clk(clk),
	.d(dffe4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_x_res_d_3),
	.prn(vcc));
defparam \cordic_x_res_d[3] .is_wysiwyg = "true";
defparam \cordic_x_res_d[3] .power_up = "low";

dffeas \cordic_x_res_2c[3] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_x_res_2c_3),
	.prn(vcc));
defparam \cordic_x_res_2c[3] .is_wysiwyg = "true";
defparam \cordic_x_res_2c[3] .power_up = "low";

dffeas \cordic_y_res_d[4] (
	.clk(clk),
	.d(pipeline_dffe_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_y_res_d_4),
	.prn(vcc));
defparam \cordic_y_res_d[4] .is_wysiwyg = "true";
defparam \cordic_y_res_d[4] .power_up = "low";

dffeas \cordic_y_res_2c[4] (
	.clk(clk),
	.d(\Add1~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_y_res_2c_4),
	.prn(vcc));
defparam \cordic_y_res_2c[4] .is_wysiwyg = "true";
defparam \cordic_y_res_2c[4] .power_up = "low";

dffeas \cordic_x_res_d[4] (
	.clk(clk),
	.d(dffe5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_x_res_d_4),
	.prn(vcc));
defparam \cordic_x_res_d[4] .is_wysiwyg = "true";
defparam \cordic_x_res_d[4] .power_up = "low";

dffeas \cordic_x_res_2c[4] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_x_res_2c_4),
	.prn(vcc));
defparam \cordic_x_res_2c[4] .is_wysiwyg = "true";
defparam \cordic_x_res_2c[4] .power_up = "low";

dffeas \cordic_y_res_d[5] (
	.clk(clk),
	.d(pipeline_dffe_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_y_res_d_5),
	.prn(vcc));
defparam \cordic_y_res_d[5] .is_wysiwyg = "true";
defparam \cordic_y_res_d[5] .power_up = "low";

dffeas \cordic_y_res_2c[5] (
	.clk(clk),
	.d(\Add1~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_y_res_2c_5),
	.prn(vcc));
defparam \cordic_y_res_2c[5] .is_wysiwyg = "true";
defparam \cordic_y_res_2c[5] .power_up = "low";

dffeas \cordic_x_res_d[5] (
	.clk(clk),
	.d(dffe6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_x_res_d_5),
	.prn(vcc));
defparam \cordic_x_res_d[5] .is_wysiwyg = "true";
defparam \cordic_x_res_d[5] .power_up = "low";

dffeas \cordic_x_res_2c[5] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_x_res_2c_5),
	.prn(vcc));
defparam \cordic_x_res_2c[5] .is_wysiwyg = "true";
defparam \cordic_x_res_2c[5] .power_up = "low";

dffeas \cordic_y_res_d[6] (
	.clk(clk),
	.d(pipeline_dffe_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_y_res_d_6),
	.prn(vcc));
defparam \cordic_y_res_d[6] .is_wysiwyg = "true";
defparam \cordic_y_res_d[6] .power_up = "low";

dffeas \cordic_y_res_2c[6] (
	.clk(clk),
	.d(\Add1~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_y_res_2c_6),
	.prn(vcc));
defparam \cordic_y_res_2c[6] .is_wysiwyg = "true";
defparam \cordic_y_res_2c[6] .power_up = "low";

dffeas \cordic_x_res_d[6] (
	.clk(clk),
	.d(dffe7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_x_res_d_6),
	.prn(vcc));
defparam \cordic_x_res_d[6] .is_wysiwyg = "true";
defparam \cordic_x_res_d[6] .power_up = "low";

dffeas \cordic_x_res_2c[6] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_x_res_2c_6),
	.prn(vcc));
defparam \cordic_x_res_2c[6] .is_wysiwyg = "true";
defparam \cordic_x_res_2c[6] .power_up = "low";

dffeas \cordic_y_res_d[7] (
	.clk(clk),
	.d(pipeline_dffe_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_y_res_d_7),
	.prn(vcc));
defparam \cordic_y_res_d[7] .is_wysiwyg = "true";
defparam \cordic_y_res_d[7] .power_up = "low";

dffeas \cordic_y_res_2c[7] (
	.clk(clk),
	.d(\Add1~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_y_res_2c_7),
	.prn(vcc));
defparam \cordic_y_res_2c[7] .is_wysiwyg = "true";
defparam \cordic_y_res_2c[7] .power_up = "low";

dffeas \cordic_x_res_d[7] (
	.clk(clk),
	.d(dffe8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_x_res_d_7),
	.prn(vcc));
defparam \cordic_x_res_d[7] .is_wysiwyg = "true";
defparam \cordic_x_res_d[7] .power_up = "low";

dffeas \cordic_x_res_2c[7] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_x_res_2c_7),
	.prn(vcc));
defparam \cordic_x_res_2c[7] .is_wysiwyg = "true";
defparam \cordic_x_res_2c[7] .power_up = "low";

dffeas \cordic_y_res_d[8] (
	.clk(clk),
	.d(pipeline_dffe_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_y_res_d_8),
	.prn(vcc));
defparam \cordic_y_res_d[8] .is_wysiwyg = "true";
defparam \cordic_y_res_d[8] .power_up = "low";

dffeas \cordic_y_res_2c[8] (
	.clk(clk),
	.d(\Add1~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_y_res_2c_8),
	.prn(vcc));
defparam \cordic_y_res_2c[8] .is_wysiwyg = "true";
defparam \cordic_y_res_2c[8] .power_up = "low";

dffeas \cordic_x_res_d[8] (
	.clk(clk),
	.d(dffe9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_x_res_d_8),
	.prn(vcc));
defparam \cordic_x_res_d[8] .is_wysiwyg = "true";
defparam \cordic_x_res_d[8] .power_up = "low";

dffeas \cordic_x_res_2c[8] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_x_res_2c_8),
	.prn(vcc));
defparam \cordic_x_res_2c[8] .is_wysiwyg = "true";
defparam \cordic_x_res_2c[8] .power_up = "low";

dffeas \cordic_y_res_d[9] (
	.clk(clk),
	.d(pipeline_dffe_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_y_res_d_9),
	.prn(vcc));
defparam \cordic_y_res_d[9] .is_wysiwyg = "true";
defparam \cordic_y_res_d[9] .power_up = "low";

dffeas \cordic_y_res_2c[9] (
	.clk(clk),
	.d(\Add1~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_y_res_2c_9),
	.prn(vcc));
defparam \cordic_y_res_2c[9] .is_wysiwyg = "true";
defparam \cordic_y_res_2c[9] .power_up = "low";

dffeas \cordic_x_res_d[9] (
	.clk(clk),
	.d(dffe10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_x_res_d_9),
	.prn(vcc));
defparam \cordic_x_res_d[9] .is_wysiwyg = "true";
defparam \cordic_x_res_d[9] .power_up = "low";

dffeas \cordic_x_res_2c[9] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_x_res_2c_9),
	.prn(vcc));
defparam \cordic_x_res_2c[9] .is_wysiwyg = "true";
defparam \cordic_x_res_2c[9] .power_up = "low";

dffeas \cordic_y_res_d[10] (
	.clk(clk),
	.d(pipeline_dffe_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_y_res_d_10),
	.prn(vcc));
defparam \cordic_y_res_d[10] .is_wysiwyg = "true";
defparam \cordic_y_res_d[10] .power_up = "low";

dffeas \cordic_y_res_2c[10] (
	.clk(clk),
	.d(\Add1~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_y_res_2c_10),
	.prn(vcc));
defparam \cordic_y_res_2c[10] .is_wysiwyg = "true";
defparam \cordic_y_res_2c[10] .power_up = "low";

dffeas \cordic_x_res_d[10] (
	.clk(clk),
	.d(dffe11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_x_res_d_10),
	.prn(vcc));
defparam \cordic_x_res_d[10] .is_wysiwyg = "true";
defparam \cordic_x_res_d[10] .power_up = "low";

dffeas \cordic_x_res_2c[10] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_x_res_2c_10),
	.prn(vcc));
defparam \cordic_x_res_2c[10] .is_wysiwyg = "true";
defparam \cordic_x_res_2c[10] .power_up = "low";

dffeas \cordic_y_res_d[11] (
	.clk(clk),
	.d(pipeline_dffe_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_y_res_d_11),
	.prn(vcc));
defparam \cordic_y_res_d[11] .is_wysiwyg = "true";
defparam \cordic_y_res_d[11] .power_up = "low";

dffeas \cordic_y_res_2c[11] (
	.clk(clk),
	.d(\Add1~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_y_res_2c_11),
	.prn(vcc));
defparam \cordic_y_res_2c[11] .is_wysiwyg = "true";
defparam \cordic_y_res_2c[11] .power_up = "low";

dffeas \cordic_x_res_d[11] (
	.clk(clk),
	.d(dffe12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_x_res_d_11),
	.prn(vcc));
defparam \cordic_x_res_d[11] .is_wysiwyg = "true";
defparam \cordic_x_res_d[11] .power_up = "low";

dffeas \cordic_x_res_2c[11] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_x_res_2c_11),
	.prn(vcc));
defparam \cordic_x_res_2c[11] .is_wysiwyg = "true";
defparam \cordic_x_res_2c[11] .power_up = "low";

dffeas \cordic_y_res_d[12] (
	.clk(clk),
	.d(pipeline_dffe_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_y_res_d_12),
	.prn(vcc));
defparam \cordic_y_res_d[12] .is_wysiwyg = "true";
defparam \cordic_y_res_d[12] .power_up = "low";

dffeas \cordic_y_res_2c[12] (
	.clk(clk),
	.d(\Add1~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_y_res_2c_12),
	.prn(vcc));
defparam \cordic_y_res_2c[12] .is_wysiwyg = "true";
defparam \cordic_y_res_2c[12] .power_up = "low";

dffeas \cordic_x_res_d[12] (
	.clk(clk),
	.d(dffe13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_x_res_d_12),
	.prn(vcc));
defparam \cordic_x_res_d[12] .is_wysiwyg = "true";
defparam \cordic_x_res_d[12] .power_up = "low";

dffeas \cordic_x_res_2c[12] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_x_res_2c_12),
	.prn(vcc));
defparam \cordic_x_res_2c[12] .is_wysiwyg = "true";
defparam \cordic_x_res_2c[12] .power_up = "low";

dffeas \cordic_y_res_d[13] (
	.clk(clk),
	.d(pipeline_dffe_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_y_res_d_13),
	.prn(vcc));
defparam \cordic_y_res_d[13] .is_wysiwyg = "true";
defparam \cordic_y_res_d[13] .power_up = "low";

dffeas \cordic_y_res_2c[13] (
	.clk(clk),
	.d(\Add1~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_y_res_2c_13),
	.prn(vcc));
defparam \cordic_y_res_2c[13] .is_wysiwyg = "true";
defparam \cordic_y_res_2c[13] .power_up = "low";

dffeas \cordic_x_res_d[13] (
	.clk(clk),
	.d(dffe14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_x_res_d_13),
	.prn(vcc));
defparam \cordic_x_res_d[13] .is_wysiwyg = "true";
defparam \cordic_x_res_d[13] .power_up = "low";

dffeas \cordic_x_res_2c[13] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_x_res_2c_13),
	.prn(vcc));
defparam \cordic_x_res_2c[13] .is_wysiwyg = "true";
defparam \cordic_x_res_2c[13] .power_up = "low";

dffeas \cordic_y_res_d[14] (
	.clk(clk),
	.d(pipeline_dffe_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_y_res_d_14),
	.prn(vcc));
defparam \cordic_y_res_d[14] .is_wysiwyg = "true";
defparam \cordic_y_res_d[14] .power_up = "low";

dffeas \cordic_y_res_2c[14] (
	.clk(clk),
	.d(\Add1~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_y_res_2c_14),
	.prn(vcc));
defparam \cordic_y_res_2c[14] .is_wysiwyg = "true";
defparam \cordic_y_res_2c[14] .power_up = "low";

dffeas \cordic_x_res_d[14] (
	.clk(clk),
	.d(dffe15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_x_res_d_14),
	.prn(vcc));
defparam \cordic_x_res_d[14] .is_wysiwyg = "true";
defparam \cordic_x_res_d[14] .power_up = "low";

dffeas \cordic_x_res_2c[14] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_x_res_2c_14),
	.prn(vcc));
defparam \cordic_x_res_2c[14] .is_wysiwyg = "true";
defparam \cordic_x_res_2c[14] .power_up = "low";

dffeas \cordic_y_res_d[15] (
	.clk(clk),
	.d(pipeline_dffe_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_y_res_d_15),
	.prn(vcc));
defparam \cordic_y_res_d[15] .is_wysiwyg = "true";
defparam \cordic_y_res_d[15] .power_up = "low";

dffeas \cordic_y_res_2c[15] (
	.clk(clk),
	.d(\Add1~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_y_res_2c_15),
	.prn(vcc));
defparam \cordic_y_res_2c[15] .is_wysiwyg = "true";
defparam \cordic_y_res_2c[15] .power_up = "low";

dffeas \cordic_x_res_d[15] (
	.clk(clk),
	.d(dffe16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_x_res_d_15),
	.prn(vcc));
defparam \cordic_x_res_d[15] .is_wysiwyg = "true";
defparam \cordic_x_res_d[15] .power_up = "low";

dffeas \cordic_x_res_2c[15] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_x_res_2c_15),
	.prn(vcc));
defparam \cordic_x_res_2c[15] .is_wysiwyg = "true";
defparam \cordic_x_res_2c[15] .power_up = "low";

dffeas \cordic_y_res_d[16] (
	.clk(clk),
	.d(pipeline_dffe_16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_y_res_d_16),
	.prn(vcc));
defparam \cordic_y_res_d[16] .is_wysiwyg = "true";
defparam \cordic_y_res_d[16] .power_up = "low";

dffeas \cordic_y_res_2c[16] (
	.clk(clk),
	.d(\Add1~65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_y_res_2c_16),
	.prn(vcc));
defparam \cordic_y_res_2c[16] .is_wysiwyg = "true";
defparam \cordic_y_res_2c[16] .power_up = "low";

dffeas \cordic_x_res_d[16] (
	.clk(clk),
	.d(dffe17),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_x_res_d_16),
	.prn(vcc));
defparam \cordic_x_res_d[16] .is_wysiwyg = "true";
defparam \cordic_x_res_d[16] .power_up = "low";

dffeas \cordic_x_res_2c[16] (
	.clk(clk),
	.d(\Add0~65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_x_res_2c_16),
	.prn(vcc));
defparam \cordic_x_res_2c[16] .is_wysiwyg = "true";
defparam \cordic_x_res_2c[16] .power_up = "low";

dffeas \cordic_y_res_d[17] (
	.clk(clk),
	.d(pipeline_dffe_17),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_y_res_d_17),
	.prn(vcc));
defparam \cordic_y_res_d[17] .is_wysiwyg = "true";
defparam \cordic_y_res_d[17] .power_up = "low";

dffeas \cordic_y_res_2c[17] (
	.clk(clk),
	.d(\Add1~69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_y_res_2c_17),
	.prn(vcc));
defparam \cordic_y_res_2c[17] .is_wysiwyg = "true";
defparam \cordic_y_res_2c[17] .power_up = "low";

dffeas \cordic_x_res_d[17] (
	.clk(clk),
	.d(dffe18),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_x_res_d_17),
	.prn(vcc));
defparam \cordic_x_res_d[17] .is_wysiwyg = "true";
defparam \cordic_x_res_d[17] .power_up = "low";

dffeas \cordic_x_res_2c[17] (
	.clk(clk),
	.d(\Add0~69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cordic_x_res_2c_17),
	.prn(vcc));
defparam \cordic_x_res_2c[17] .is_wysiwyg = "true";
defparam \cordic_x_res_2c[17] .power_up = "low";

arriav_lcell_comb \Add1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~1_sumout ),
	.cout(\Add1~2 ),
	.shareout());
defparam \Add1~1 .extended_lut = "off";
defparam \Add1~1 .lut_mask = 64'h000000000000FF00;
defparam \Add1~1 .shared_arith = "off";

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "off";

arriav_lcell_comb \Add1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~5_sumout ),
	.cout(\Add1~6 ),
	.shareout());
defparam \Add1~5 .extended_lut = "off";
defparam \Add1~5 .lut_mask = 64'h000000000000FF00;
defparam \Add1~5 .shared_arith = "off";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000000000FF00;
defparam \Add0~5 .shared_arith = "off";

arriav_lcell_comb \Add1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~9_sumout ),
	.cout(\Add1~10 ),
	.shareout());
defparam \Add1~9 .extended_lut = "off";
defparam \Add1~9 .lut_mask = 64'h000000000000FF00;
defparam \Add1~9 .shared_arith = "off";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000000000FF00;
defparam \Add0~9 .shared_arith = "off";

arriav_lcell_comb \Add1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~13_sumout ),
	.cout(\Add1~14 ),
	.shareout());
defparam \Add1~13 .extended_lut = "off";
defparam \Add1~13 .lut_mask = 64'h000000000000FF00;
defparam \Add1~13 .shared_arith = "off";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000000000FF00;
defparam \Add0~13 .shared_arith = "off";

arriav_lcell_comb \Add1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~17_sumout ),
	.cout(\Add1~18 ),
	.shareout());
defparam \Add1~17 .extended_lut = "off";
defparam \Add1~17 .lut_mask = 64'h000000000000FF00;
defparam \Add1~17 .shared_arith = "off";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000000000FF00;
defparam \Add0~17 .shared_arith = "off";

arriav_lcell_comb \Add1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~21_sumout ),
	.cout(\Add1~22 ),
	.shareout());
defparam \Add1~21 .extended_lut = "off";
defparam \Add1~21 .lut_mask = 64'h000000000000FF00;
defparam \Add1~21 .shared_arith = "off";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000000000FF00;
defparam \Add0~21 .shared_arith = "off";

arriav_lcell_comb \Add1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~25_sumout ),
	.cout(\Add1~26 ),
	.shareout());
defparam \Add1~25 .extended_lut = "off";
defparam \Add1~25 .lut_mask = 64'h000000000000FF00;
defparam \Add1~25 .shared_arith = "off";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000000000FF00;
defparam \Add0~25 .shared_arith = "off";

arriav_lcell_comb \Add1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~29_sumout ),
	.cout(\Add1~30 ),
	.shareout());
defparam \Add1~29 .extended_lut = "off";
defparam \Add1~29 .lut_mask = 64'h000000000000FF00;
defparam \Add1~29 .shared_arith = "off";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000000000FF00;
defparam \Add0~29 .shared_arith = "off";

arriav_lcell_comb \Add1~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~33_sumout ),
	.cout(\Add1~34 ),
	.shareout());
defparam \Add1~33 .extended_lut = "off";
defparam \Add1~33 .lut_mask = 64'h000000000000FF00;
defparam \Add1~33 .shared_arith = "off";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h000000000000FF00;
defparam \Add0~33 .shared_arith = "off";

arriav_lcell_comb \Add1~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~37_sumout ),
	.cout(\Add1~38 ),
	.shareout());
defparam \Add1~37 .extended_lut = "off";
defparam \Add1~37 .lut_mask = 64'h000000000000FF00;
defparam \Add1~37 .shared_arith = "off";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000000000FF00;
defparam \Add0~37 .shared_arith = "off";

arriav_lcell_comb \Add1~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~41_sumout ),
	.cout(\Add1~42 ),
	.shareout());
defparam \Add1~41 .extended_lut = "off";
defparam \Add1~41 .lut_mask = 64'h000000000000FF00;
defparam \Add1~41 .shared_arith = "off";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000000000FF00;
defparam \Add0~41 .shared_arith = "off";

arriav_lcell_comb \Add1~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~45_sumout ),
	.cout(\Add1~46 ),
	.shareout());
defparam \Add1~45 .extended_lut = "off";
defparam \Add1~45 .lut_mask = 64'h000000000000FF00;
defparam \Add1~45 .shared_arith = "off";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000000000FF00;
defparam \Add0~45 .shared_arith = "off";

arriav_lcell_comb \Add1~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~49_sumout ),
	.cout(\Add1~50 ),
	.shareout());
defparam \Add1~49 .extended_lut = "off";
defparam \Add1~49 .lut_mask = 64'h000000000000FF00;
defparam \Add1~49 .shared_arith = "off";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout());
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h000000000000FF00;
defparam \Add0~49 .shared_arith = "off";

arriav_lcell_comb \Add1~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~53_sumout ),
	.cout(\Add1~54 ),
	.shareout());
defparam \Add1~53 .extended_lut = "off";
defparam \Add1~53 .lut_mask = 64'h000000000000FF00;
defparam \Add1~53 .shared_arith = "off";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe14),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout());
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h000000000000FF00;
defparam \Add0~53 .shared_arith = "off";

arriav_lcell_comb \Add1~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_14),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~57_sumout ),
	.cout(\Add1~58 ),
	.shareout());
defparam \Add1~57 .extended_lut = "off";
defparam \Add1~57 .lut_mask = 64'h000000000000FF00;
defparam \Add1~57 .shared_arith = "off";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe15),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout());
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h000000000000FF00;
defparam \Add0~57 .shared_arith = "off";

arriav_lcell_comb \Add1~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_15),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~61_sumout ),
	.cout(\Add1~62 ),
	.shareout());
defparam \Add1~61 .extended_lut = "off";
defparam \Add1~61 .lut_mask = 64'h000000000000FF00;
defparam \Add1~61 .shared_arith = "off";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe16),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout());
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h000000000000FF00;
defparam \Add0~61 .shared_arith = "off";

arriav_lcell_comb \Add1~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_16),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~65_sumout ),
	.cout(\Add1~66 ),
	.shareout());
defparam \Add1~65 .extended_lut = "off";
defparam \Add1~65 .lut_mask = 64'h000000000000FF00;
defparam \Add1~65 .shared_arith = "off";

arriav_lcell_comb \Add0~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe17),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~65_sumout ),
	.cout(\Add0~66 ),
	.shareout());
defparam \Add0~65 .extended_lut = "off";
defparam \Add0~65 .lut_mask = 64'h000000000000FF00;
defparam \Add0~65 .shared_arith = "off";

arriav_lcell_comb \Add1~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_17),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add1~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add1~69_sumout ),
	.cout(),
	.shareout());
defparam \Add1~69 .extended_lut = "off";
defparam \Add1~69 .lut_mask = 64'h000000000000FF00;
defparam \Add1~69 .shared_arith = "off";

arriav_lcell_comb \Add0~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe18),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~69_sumout ),
	.cout(),
	.shareout());
defparam \Add0~69 .extended_lut = "off";
defparam \Add0~69 .lut_mask = 64'h000000000000FF00;
defparam \Add0~69 .shared_arith = "off";

endmodule

module nco_test_cord_fs (
	cor1x_10,
	sin_o_0,
	corx_10,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	cor1x_10;
input 	sin_o_0;
input 	corx_10;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \cor1x[10] (
	.clk(clk),
	.d(corx_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(cor1x_10),
	.prn(vcc));
defparam \cor1x[10] .is_wysiwyg = "true";
defparam \cor1x[10] .power_up = "low";

endmodule

module nco_test_cord_init (
	corz_14,
	dxxpdo_18,
	corz_13,
	dxxpdo_17,
	corz_12,
	dxxpdo_16,
	corz_11,
	dxxpdo_15,
	corz_10,
	dxxpdo_14,
	corz_9,
	dxxpdo_13,
	corz_8,
	dxxpdo_12,
	corz_7,
	dxxpdo_11,
	corz_6,
	dxxpdo_10,
	corz_5,
	dxxpdo_9,
	corz_4,
	dxxpdo_8,
	corz_3,
	dxxpdo_7,
	corz_2,
	dxxpdo_6,
	corz_1,
	dxxpdo_5,
	corz_0,
	dxxpdo_4,
	sin_o_0,
	corx_10,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	corz_14;
input 	dxxpdo_18;
output 	corz_13;
input 	dxxpdo_17;
output 	corz_12;
input 	dxxpdo_16;
output 	corz_11;
input 	dxxpdo_15;
output 	corz_10;
input 	dxxpdo_14;
output 	corz_9;
input 	dxxpdo_13;
output 	corz_8;
input 	dxxpdo_12;
output 	corz_7;
input 	dxxpdo_11;
output 	corz_6;
input 	dxxpdo_10;
output 	corz_5;
input 	dxxpdo_9;
output 	corz_4;
input 	dxxpdo_8;
output 	corz_3;
input 	dxxpdo_7;
output 	corz_2;
input 	dxxpdo_6;
output 	corz_1;
input 	dxxpdo_5;
output 	corz_0;
input 	dxxpdo_4;
input 	sin_o_0;
output 	corx_10;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \corx[10]~0_combout ;


dffeas \corz[14] (
	.clk(clk),
	.d(dxxpdo_18),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(corz_14),
	.prn(vcc));
defparam \corz[14] .is_wysiwyg = "true";
defparam \corz[14] .power_up = "low";

dffeas \corz[13] (
	.clk(clk),
	.d(dxxpdo_17),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(corz_13),
	.prn(vcc));
defparam \corz[13] .is_wysiwyg = "true";
defparam \corz[13] .power_up = "low";

dffeas \corz[12] (
	.clk(clk),
	.d(dxxpdo_16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(corz_12),
	.prn(vcc));
defparam \corz[12] .is_wysiwyg = "true";
defparam \corz[12] .power_up = "low";

dffeas \corz[11] (
	.clk(clk),
	.d(dxxpdo_15),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(corz_11),
	.prn(vcc));
defparam \corz[11] .is_wysiwyg = "true";
defparam \corz[11] .power_up = "low";

dffeas \corz[10] (
	.clk(clk),
	.d(dxxpdo_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(corz_10),
	.prn(vcc));
defparam \corz[10] .is_wysiwyg = "true";
defparam \corz[10] .power_up = "low";

dffeas \corz[9] (
	.clk(clk),
	.d(dxxpdo_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(corz_9),
	.prn(vcc));
defparam \corz[9] .is_wysiwyg = "true";
defparam \corz[9] .power_up = "low";

dffeas \corz[8] (
	.clk(clk),
	.d(dxxpdo_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(corz_8),
	.prn(vcc));
defparam \corz[8] .is_wysiwyg = "true";
defparam \corz[8] .power_up = "low";

dffeas \corz[7] (
	.clk(clk),
	.d(dxxpdo_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(corz_7),
	.prn(vcc));
defparam \corz[7] .is_wysiwyg = "true";
defparam \corz[7] .power_up = "low";

dffeas \corz[6] (
	.clk(clk),
	.d(dxxpdo_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(corz_6),
	.prn(vcc));
defparam \corz[6] .is_wysiwyg = "true";
defparam \corz[6] .power_up = "low";

dffeas \corz[5] (
	.clk(clk),
	.d(dxxpdo_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(corz_5),
	.prn(vcc));
defparam \corz[5] .is_wysiwyg = "true";
defparam \corz[5] .power_up = "low";

dffeas \corz[4] (
	.clk(clk),
	.d(dxxpdo_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(corz_4),
	.prn(vcc));
defparam \corz[4] .is_wysiwyg = "true";
defparam \corz[4] .power_up = "low";

dffeas \corz[3] (
	.clk(clk),
	.d(dxxpdo_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(corz_3),
	.prn(vcc));
defparam \corz[3] .is_wysiwyg = "true";
defparam \corz[3] .power_up = "low";

dffeas \corz[2] (
	.clk(clk),
	.d(dxxpdo_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(corz_2),
	.prn(vcc));
defparam \corz[2] .is_wysiwyg = "true";
defparam \corz[2] .power_up = "low";

dffeas \corz[1] (
	.clk(clk),
	.d(dxxpdo_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(corz_1),
	.prn(vcc));
defparam \corz[1] .is_wysiwyg = "true";
defparam \corz[1] .power_up = "low";

dffeas \corz[0] (
	.clk(clk),
	.d(dxxpdo_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(corz_0),
	.prn(vcc));
defparam \corz[0] .is_wysiwyg = "true";
defparam \corz[0] .power_up = "low";

dffeas \corx[10] (
	.clk(clk),
	.d(\corx[10]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(corx_10),
	.prn(vcc));
defparam \corx[10] .is_wysiwyg = "true";
defparam \corx[10] .power_up = "low";

arriav_lcell_comb \corx[10]~0 (
	.dataa(!reset_n),
	.datab(!clken),
	.datac(!corx_10),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\corx[10]~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \corx[10]~0 .extended_lut = "off";
defparam \corx[10]~0 .lut_mask = 64'h7F7F7F7F7F7F7F7F;
defparam \corx[10]~0 .shared_arith = "off";

endmodule

module nco_test_cord_seg_sel (
	seg_rot_1,
	seg_rot_0,
	dxxpdo_20,
	dxxpdo_19,
	sin_o_0,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	seg_rot_1;
output 	seg_rot_0;
input 	dxxpdo_20;
input 	dxxpdo_19;
input 	sin_o_0;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \zheld[0][1]~q ;
wire \zheld[1][1]~q ;
wire \zheld[2][1]~q ;
wire \zheld[3][1]~q ;
wire \zheld[4][1]~q ;
wire \zheld[5][1]~q ;
wire \zheld[6][1]~q ;
wire \zheld[7][1]~q ;
wire \zheld[8][1]~q ;
wire \zheld[9][1]~q ;
wire \zheld[10][1]~q ;
wire \zheld[11][1]~q ;
wire \zheld[12][1]~q ;
wire \zheld[13][1]~q ;
wire \zheld[14][1]~q ;
wire \zheld[15][1]~q ;
wire \zheld[16][1]~q ;
wire \zheld[17][1]~q ;
wire \zheld[18][1]~q ;
wire \zheld[19][1]~q ;
wire \zheld[20][1]~q ;
wire \zheld[21][1]~q ;
wire \zheld[22][1]~q ;
wire \zheld[23][1]~q ;
wire \zheld[24][1]~q ;
wire \zheld[25][1]~q ;
wire \zheld[26][1]~q ;
wire \zheld[27][1]~q ;
wire \zheld[28][1]~q ;
wire \zheld[29][1]~q ;
wire \zheld[30][1]~q ;
wire \zheld[31][1]~q ;
wire \zheld[32][1]~q ;
wire \zheld[33][1]~q ;
wire \zheld[34][1]~q ;
wire \zheld[35][1]~q ;
wire \zheld[36][1]~q ;
wire \zheld[0][0]~q ;
wire \zheld[1][0]~q ;
wire \zheld[2][0]~q ;
wire \zheld[3][0]~q ;
wire \zheld[4][0]~q ;
wire \zheld[5][0]~q ;
wire \zheld[6][0]~q ;
wire \zheld[7][0]~q ;
wire \zheld[8][0]~q ;
wire \zheld[9][0]~q ;
wire \zheld[10][0]~q ;
wire \zheld[11][0]~q ;
wire \zheld[12][0]~q ;
wire \zheld[13][0]~q ;
wire \zheld[14][0]~q ;
wire \zheld[15][0]~q ;
wire \zheld[16][0]~q ;
wire \zheld[17][0]~q ;
wire \zheld[18][0]~q ;
wire \zheld[19][0]~q ;
wire \zheld[20][0]~q ;
wire \zheld[21][0]~q ;
wire \zheld[22][0]~q ;
wire \zheld[23][0]~q ;
wire \zheld[24][0]~q ;
wire \zheld[25][0]~q ;
wire \zheld[26][0]~q ;
wire \zheld[27][0]~q ;
wire \zheld[28][0]~q ;
wire \zheld[29][0]~q ;
wire \zheld[30][0]~q ;
wire \zheld[31][0]~q ;
wire \zheld[32][0]~q ;
wire \zheld[33][0]~q ;
wire \zheld[34][0]~q ;
wire \zheld[35][0]~q ;
wire \zheld[36][0]~q ;


dffeas \seg_rot[1] (
	.clk(clk),
	.d(\zheld[36][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(seg_rot_1),
	.prn(vcc));
defparam \seg_rot[1] .is_wysiwyg = "true";
defparam \seg_rot[1] .power_up = "low";

dffeas \seg_rot[0] (
	.clk(clk),
	.d(\zheld[36][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(seg_rot_0),
	.prn(vcc));
defparam \seg_rot[0] .is_wysiwyg = "true";
defparam \seg_rot[0] .power_up = "low";

dffeas \zheld[0][1] (
	.clk(clk),
	.d(dxxpdo_20),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[0][1]~q ),
	.prn(vcc));
defparam \zheld[0][1] .is_wysiwyg = "true";
defparam \zheld[0][1] .power_up = "low";

dffeas \zheld[1][1] (
	.clk(clk),
	.d(\zheld[0][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[1][1]~q ),
	.prn(vcc));
defparam \zheld[1][1] .is_wysiwyg = "true";
defparam \zheld[1][1] .power_up = "low";

dffeas \zheld[2][1] (
	.clk(clk),
	.d(\zheld[1][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[2][1]~q ),
	.prn(vcc));
defparam \zheld[2][1] .is_wysiwyg = "true";
defparam \zheld[2][1] .power_up = "low";

dffeas \zheld[3][1] (
	.clk(clk),
	.d(\zheld[2][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[3][1]~q ),
	.prn(vcc));
defparam \zheld[3][1] .is_wysiwyg = "true";
defparam \zheld[3][1] .power_up = "low";

dffeas \zheld[4][1] (
	.clk(clk),
	.d(\zheld[3][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[4][1]~q ),
	.prn(vcc));
defparam \zheld[4][1] .is_wysiwyg = "true";
defparam \zheld[4][1] .power_up = "low";

dffeas \zheld[5][1] (
	.clk(clk),
	.d(\zheld[4][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[5][1]~q ),
	.prn(vcc));
defparam \zheld[5][1] .is_wysiwyg = "true";
defparam \zheld[5][1] .power_up = "low";

dffeas \zheld[6][1] (
	.clk(clk),
	.d(\zheld[5][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[6][1]~q ),
	.prn(vcc));
defparam \zheld[6][1] .is_wysiwyg = "true";
defparam \zheld[6][1] .power_up = "low";

dffeas \zheld[7][1] (
	.clk(clk),
	.d(\zheld[6][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[7][1]~q ),
	.prn(vcc));
defparam \zheld[7][1] .is_wysiwyg = "true";
defparam \zheld[7][1] .power_up = "low";

dffeas \zheld[8][1] (
	.clk(clk),
	.d(\zheld[7][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[8][1]~q ),
	.prn(vcc));
defparam \zheld[8][1] .is_wysiwyg = "true";
defparam \zheld[8][1] .power_up = "low";

dffeas \zheld[9][1] (
	.clk(clk),
	.d(\zheld[8][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[9][1]~q ),
	.prn(vcc));
defparam \zheld[9][1] .is_wysiwyg = "true";
defparam \zheld[9][1] .power_up = "low";

dffeas \zheld[10][1] (
	.clk(clk),
	.d(\zheld[9][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[10][1]~q ),
	.prn(vcc));
defparam \zheld[10][1] .is_wysiwyg = "true";
defparam \zheld[10][1] .power_up = "low";

dffeas \zheld[11][1] (
	.clk(clk),
	.d(\zheld[10][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[11][1]~q ),
	.prn(vcc));
defparam \zheld[11][1] .is_wysiwyg = "true";
defparam \zheld[11][1] .power_up = "low";

dffeas \zheld[12][1] (
	.clk(clk),
	.d(\zheld[11][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[12][1]~q ),
	.prn(vcc));
defparam \zheld[12][1] .is_wysiwyg = "true";
defparam \zheld[12][1] .power_up = "low";

dffeas \zheld[13][1] (
	.clk(clk),
	.d(\zheld[12][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[13][1]~q ),
	.prn(vcc));
defparam \zheld[13][1] .is_wysiwyg = "true";
defparam \zheld[13][1] .power_up = "low";

dffeas \zheld[14][1] (
	.clk(clk),
	.d(\zheld[13][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[14][1]~q ),
	.prn(vcc));
defparam \zheld[14][1] .is_wysiwyg = "true";
defparam \zheld[14][1] .power_up = "low";

dffeas \zheld[15][1] (
	.clk(clk),
	.d(\zheld[14][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[15][1]~q ),
	.prn(vcc));
defparam \zheld[15][1] .is_wysiwyg = "true";
defparam \zheld[15][1] .power_up = "low";

dffeas \zheld[16][1] (
	.clk(clk),
	.d(\zheld[15][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[16][1]~q ),
	.prn(vcc));
defparam \zheld[16][1] .is_wysiwyg = "true";
defparam \zheld[16][1] .power_up = "low";

dffeas \zheld[17][1] (
	.clk(clk),
	.d(\zheld[16][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[17][1]~q ),
	.prn(vcc));
defparam \zheld[17][1] .is_wysiwyg = "true";
defparam \zheld[17][1] .power_up = "low";

dffeas \zheld[18][1] (
	.clk(clk),
	.d(\zheld[17][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[18][1]~q ),
	.prn(vcc));
defparam \zheld[18][1] .is_wysiwyg = "true";
defparam \zheld[18][1] .power_up = "low";

dffeas \zheld[19][1] (
	.clk(clk),
	.d(\zheld[18][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[19][1]~q ),
	.prn(vcc));
defparam \zheld[19][1] .is_wysiwyg = "true";
defparam \zheld[19][1] .power_up = "low";

dffeas \zheld[20][1] (
	.clk(clk),
	.d(\zheld[19][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[20][1]~q ),
	.prn(vcc));
defparam \zheld[20][1] .is_wysiwyg = "true";
defparam \zheld[20][1] .power_up = "low";

dffeas \zheld[21][1] (
	.clk(clk),
	.d(\zheld[20][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[21][1]~q ),
	.prn(vcc));
defparam \zheld[21][1] .is_wysiwyg = "true";
defparam \zheld[21][1] .power_up = "low";

dffeas \zheld[22][1] (
	.clk(clk),
	.d(\zheld[21][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[22][1]~q ),
	.prn(vcc));
defparam \zheld[22][1] .is_wysiwyg = "true";
defparam \zheld[22][1] .power_up = "low";

dffeas \zheld[23][1] (
	.clk(clk),
	.d(\zheld[22][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[23][1]~q ),
	.prn(vcc));
defparam \zheld[23][1] .is_wysiwyg = "true";
defparam \zheld[23][1] .power_up = "low";

dffeas \zheld[24][1] (
	.clk(clk),
	.d(\zheld[23][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[24][1]~q ),
	.prn(vcc));
defparam \zheld[24][1] .is_wysiwyg = "true";
defparam \zheld[24][1] .power_up = "low";

dffeas \zheld[25][1] (
	.clk(clk),
	.d(\zheld[24][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[25][1]~q ),
	.prn(vcc));
defparam \zheld[25][1] .is_wysiwyg = "true";
defparam \zheld[25][1] .power_up = "low";

dffeas \zheld[26][1] (
	.clk(clk),
	.d(\zheld[25][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[26][1]~q ),
	.prn(vcc));
defparam \zheld[26][1] .is_wysiwyg = "true";
defparam \zheld[26][1] .power_up = "low";

dffeas \zheld[27][1] (
	.clk(clk),
	.d(\zheld[26][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[27][1]~q ),
	.prn(vcc));
defparam \zheld[27][1] .is_wysiwyg = "true";
defparam \zheld[27][1] .power_up = "low";

dffeas \zheld[28][1] (
	.clk(clk),
	.d(\zheld[27][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[28][1]~q ),
	.prn(vcc));
defparam \zheld[28][1] .is_wysiwyg = "true";
defparam \zheld[28][1] .power_up = "low";

dffeas \zheld[29][1] (
	.clk(clk),
	.d(\zheld[28][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[29][1]~q ),
	.prn(vcc));
defparam \zheld[29][1] .is_wysiwyg = "true";
defparam \zheld[29][1] .power_up = "low";

dffeas \zheld[30][1] (
	.clk(clk),
	.d(\zheld[29][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[30][1]~q ),
	.prn(vcc));
defparam \zheld[30][1] .is_wysiwyg = "true";
defparam \zheld[30][1] .power_up = "low";

dffeas \zheld[31][1] (
	.clk(clk),
	.d(\zheld[30][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[31][1]~q ),
	.prn(vcc));
defparam \zheld[31][1] .is_wysiwyg = "true";
defparam \zheld[31][1] .power_up = "low";

dffeas \zheld[32][1] (
	.clk(clk),
	.d(\zheld[31][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[32][1]~q ),
	.prn(vcc));
defparam \zheld[32][1] .is_wysiwyg = "true";
defparam \zheld[32][1] .power_up = "low";

dffeas \zheld[33][1] (
	.clk(clk),
	.d(\zheld[32][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[33][1]~q ),
	.prn(vcc));
defparam \zheld[33][1] .is_wysiwyg = "true";
defparam \zheld[33][1] .power_up = "low";

dffeas \zheld[34][1] (
	.clk(clk),
	.d(\zheld[33][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[34][1]~q ),
	.prn(vcc));
defparam \zheld[34][1] .is_wysiwyg = "true";
defparam \zheld[34][1] .power_up = "low";

dffeas \zheld[35][1] (
	.clk(clk),
	.d(\zheld[34][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[35][1]~q ),
	.prn(vcc));
defparam \zheld[35][1] .is_wysiwyg = "true";
defparam \zheld[35][1] .power_up = "low";

dffeas \zheld[36][1] (
	.clk(clk),
	.d(\zheld[35][1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[36][1]~q ),
	.prn(vcc));
defparam \zheld[36][1] .is_wysiwyg = "true";
defparam \zheld[36][1] .power_up = "low";

dffeas \zheld[0][0] (
	.clk(clk),
	.d(dxxpdo_19),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[0][0]~q ),
	.prn(vcc));
defparam \zheld[0][0] .is_wysiwyg = "true";
defparam \zheld[0][0] .power_up = "low";

dffeas \zheld[1][0] (
	.clk(clk),
	.d(\zheld[0][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[1][0]~q ),
	.prn(vcc));
defparam \zheld[1][0] .is_wysiwyg = "true";
defparam \zheld[1][0] .power_up = "low";

dffeas \zheld[2][0] (
	.clk(clk),
	.d(\zheld[1][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[2][0]~q ),
	.prn(vcc));
defparam \zheld[2][0] .is_wysiwyg = "true";
defparam \zheld[2][0] .power_up = "low";

dffeas \zheld[3][0] (
	.clk(clk),
	.d(\zheld[2][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[3][0]~q ),
	.prn(vcc));
defparam \zheld[3][0] .is_wysiwyg = "true";
defparam \zheld[3][0] .power_up = "low";

dffeas \zheld[4][0] (
	.clk(clk),
	.d(\zheld[3][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[4][0]~q ),
	.prn(vcc));
defparam \zheld[4][0] .is_wysiwyg = "true";
defparam \zheld[4][0] .power_up = "low";

dffeas \zheld[5][0] (
	.clk(clk),
	.d(\zheld[4][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[5][0]~q ),
	.prn(vcc));
defparam \zheld[5][0] .is_wysiwyg = "true";
defparam \zheld[5][0] .power_up = "low";

dffeas \zheld[6][0] (
	.clk(clk),
	.d(\zheld[5][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[6][0]~q ),
	.prn(vcc));
defparam \zheld[6][0] .is_wysiwyg = "true";
defparam \zheld[6][0] .power_up = "low";

dffeas \zheld[7][0] (
	.clk(clk),
	.d(\zheld[6][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[7][0]~q ),
	.prn(vcc));
defparam \zheld[7][0] .is_wysiwyg = "true";
defparam \zheld[7][0] .power_up = "low";

dffeas \zheld[8][0] (
	.clk(clk),
	.d(\zheld[7][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[8][0]~q ),
	.prn(vcc));
defparam \zheld[8][0] .is_wysiwyg = "true";
defparam \zheld[8][0] .power_up = "low";

dffeas \zheld[9][0] (
	.clk(clk),
	.d(\zheld[8][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[9][0]~q ),
	.prn(vcc));
defparam \zheld[9][0] .is_wysiwyg = "true";
defparam \zheld[9][0] .power_up = "low";

dffeas \zheld[10][0] (
	.clk(clk),
	.d(\zheld[9][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[10][0]~q ),
	.prn(vcc));
defparam \zheld[10][0] .is_wysiwyg = "true";
defparam \zheld[10][0] .power_up = "low";

dffeas \zheld[11][0] (
	.clk(clk),
	.d(\zheld[10][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[11][0]~q ),
	.prn(vcc));
defparam \zheld[11][0] .is_wysiwyg = "true";
defparam \zheld[11][0] .power_up = "low";

dffeas \zheld[12][0] (
	.clk(clk),
	.d(\zheld[11][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[12][0]~q ),
	.prn(vcc));
defparam \zheld[12][0] .is_wysiwyg = "true";
defparam \zheld[12][0] .power_up = "low";

dffeas \zheld[13][0] (
	.clk(clk),
	.d(\zheld[12][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[13][0]~q ),
	.prn(vcc));
defparam \zheld[13][0] .is_wysiwyg = "true";
defparam \zheld[13][0] .power_up = "low";

dffeas \zheld[14][0] (
	.clk(clk),
	.d(\zheld[13][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[14][0]~q ),
	.prn(vcc));
defparam \zheld[14][0] .is_wysiwyg = "true";
defparam \zheld[14][0] .power_up = "low";

dffeas \zheld[15][0] (
	.clk(clk),
	.d(\zheld[14][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[15][0]~q ),
	.prn(vcc));
defparam \zheld[15][0] .is_wysiwyg = "true";
defparam \zheld[15][0] .power_up = "low";

dffeas \zheld[16][0] (
	.clk(clk),
	.d(\zheld[15][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[16][0]~q ),
	.prn(vcc));
defparam \zheld[16][0] .is_wysiwyg = "true";
defparam \zheld[16][0] .power_up = "low";

dffeas \zheld[17][0] (
	.clk(clk),
	.d(\zheld[16][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[17][0]~q ),
	.prn(vcc));
defparam \zheld[17][0] .is_wysiwyg = "true";
defparam \zheld[17][0] .power_up = "low";

dffeas \zheld[18][0] (
	.clk(clk),
	.d(\zheld[17][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[18][0]~q ),
	.prn(vcc));
defparam \zheld[18][0] .is_wysiwyg = "true";
defparam \zheld[18][0] .power_up = "low";

dffeas \zheld[19][0] (
	.clk(clk),
	.d(\zheld[18][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[19][0]~q ),
	.prn(vcc));
defparam \zheld[19][0] .is_wysiwyg = "true";
defparam \zheld[19][0] .power_up = "low";

dffeas \zheld[20][0] (
	.clk(clk),
	.d(\zheld[19][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[20][0]~q ),
	.prn(vcc));
defparam \zheld[20][0] .is_wysiwyg = "true";
defparam \zheld[20][0] .power_up = "low";

dffeas \zheld[21][0] (
	.clk(clk),
	.d(\zheld[20][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[21][0]~q ),
	.prn(vcc));
defparam \zheld[21][0] .is_wysiwyg = "true";
defparam \zheld[21][0] .power_up = "low";

dffeas \zheld[22][0] (
	.clk(clk),
	.d(\zheld[21][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[22][0]~q ),
	.prn(vcc));
defparam \zheld[22][0] .is_wysiwyg = "true";
defparam \zheld[22][0] .power_up = "low";

dffeas \zheld[23][0] (
	.clk(clk),
	.d(\zheld[22][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[23][0]~q ),
	.prn(vcc));
defparam \zheld[23][0] .is_wysiwyg = "true";
defparam \zheld[23][0] .power_up = "low";

dffeas \zheld[24][0] (
	.clk(clk),
	.d(\zheld[23][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[24][0]~q ),
	.prn(vcc));
defparam \zheld[24][0] .is_wysiwyg = "true";
defparam \zheld[24][0] .power_up = "low";

dffeas \zheld[25][0] (
	.clk(clk),
	.d(\zheld[24][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[25][0]~q ),
	.prn(vcc));
defparam \zheld[25][0] .is_wysiwyg = "true";
defparam \zheld[25][0] .power_up = "low";

dffeas \zheld[26][0] (
	.clk(clk),
	.d(\zheld[25][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[26][0]~q ),
	.prn(vcc));
defparam \zheld[26][0] .is_wysiwyg = "true";
defparam \zheld[26][0] .power_up = "low";

dffeas \zheld[27][0] (
	.clk(clk),
	.d(\zheld[26][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[27][0]~q ),
	.prn(vcc));
defparam \zheld[27][0] .is_wysiwyg = "true";
defparam \zheld[27][0] .power_up = "low";

dffeas \zheld[28][0] (
	.clk(clk),
	.d(\zheld[27][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[28][0]~q ),
	.prn(vcc));
defparam \zheld[28][0] .is_wysiwyg = "true";
defparam \zheld[28][0] .power_up = "low";

dffeas \zheld[29][0] (
	.clk(clk),
	.d(\zheld[28][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[29][0]~q ),
	.prn(vcc));
defparam \zheld[29][0] .is_wysiwyg = "true";
defparam \zheld[29][0] .power_up = "low";

dffeas \zheld[30][0] (
	.clk(clk),
	.d(\zheld[29][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[30][0]~q ),
	.prn(vcc));
defparam \zheld[30][0] .is_wysiwyg = "true";
defparam \zheld[30][0] .power_up = "low";

dffeas \zheld[31][0] (
	.clk(clk),
	.d(\zheld[30][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[31][0]~q ),
	.prn(vcc));
defparam \zheld[31][0] .is_wysiwyg = "true";
defparam \zheld[31][0] .power_up = "low";

dffeas \zheld[32][0] (
	.clk(clk),
	.d(\zheld[31][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[32][0]~q ),
	.prn(vcc));
defparam \zheld[32][0] .is_wysiwyg = "true";
defparam \zheld[32][0] .power_up = "low";

dffeas \zheld[33][0] (
	.clk(clk),
	.d(\zheld[32][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[33][0]~q ),
	.prn(vcc));
defparam \zheld[33][0] .is_wysiwyg = "true";
defparam \zheld[33][0] .power_up = "low";

dffeas \zheld[34][0] (
	.clk(clk),
	.d(\zheld[33][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[34][0]~q ),
	.prn(vcc));
defparam \zheld[34][0] .is_wysiwyg = "true";
defparam \zheld[34][0] .power_up = "low";

dffeas \zheld[35][0] (
	.clk(clk),
	.d(\zheld[34][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[35][0]~q ),
	.prn(vcc));
defparam \zheld[35][0] .is_wysiwyg = "true";
defparam \zheld[35][0] .power_up = "low";

dffeas \zheld[36][0] (
	.clk(clk),
	.d(\zheld[35][0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\zheld[36][0]~q ),
	.prn(vcc));
defparam \zheld[36][0] .is_wysiwyg = "true";
defparam \zheld[36][0] .power_up = "low";

endmodule

module nco_test_cordic_axor_1p_lpm (
	sin_o_0,
	pipeline_dffe_17,
	pipeline_dffe_16,
	dffe16,
	dffe18,
	pipeline_dffe_15,
	pipeline_dffe_171,
	pipeline_dffe_14,
	pipeline_dffe_161,
	pipeline_dffe_13,
	dffe17,
	pipeline_dffe_151,
	pipeline_dffe_12,
	dffe161,
	pipeline_dffe_141,
	pipeline_dffe_11,
	dffe15,
	pipeline_dffe_131,
	pipeline_dffe_10,
	dffe14,
	pipeline_dffe_121,
	pipeline_dffe_9,
	dffe13,
	pipeline_dffe_111,
	pipeline_dffe_8,
	dffe12,
	pipeline_dffe_101,
	pipeline_dffe_7,
	dffe11,
	pipeline_dffe_91,
	pipeline_dffe_6,
	dffe10,
	pipeline_dffe_81,
	pipeline_dffe_4,
	pipeline_dffe_5,
	dffe9,
	pipeline_dffe_0,
	pipeline_dffe_71,
	dffe8,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_61,
	dffe7,
	pipeline_dffe_51,
	dffe6,
	dffe4,
	dffe5,
	pipeline_dffe_41,
	pipeline_dffe_31,
	pipeline_dffe_01,
	pipeline_dffe_18,
	pipeline_dffe_21,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	sin_o_0;
output 	pipeline_dffe_17;
output 	pipeline_dffe_16;
input 	dffe16;
input 	dffe18;
output 	pipeline_dffe_15;
input 	pipeline_dffe_171;
output 	pipeline_dffe_14;
input 	pipeline_dffe_161;
output 	pipeline_dffe_13;
input 	dffe17;
input 	pipeline_dffe_151;
output 	pipeline_dffe_12;
input 	dffe161;
input 	pipeline_dffe_141;
output 	pipeline_dffe_11;
input 	dffe15;
input 	pipeline_dffe_131;
output 	pipeline_dffe_10;
input 	dffe14;
input 	pipeline_dffe_121;
output 	pipeline_dffe_9;
input 	dffe13;
input 	pipeline_dffe_111;
output 	pipeline_dffe_8;
input 	dffe12;
input 	pipeline_dffe_101;
output 	pipeline_dffe_7;
input 	dffe11;
input 	pipeline_dffe_91;
output 	pipeline_dffe_6;
input 	dffe10;
input 	pipeline_dffe_81;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
input 	dffe9;
output 	pipeline_dffe_0;
input 	pipeline_dffe_71;
input 	dffe8;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
input 	pipeline_dffe_61;
input 	dffe7;
input 	pipeline_dffe_51;
input 	dffe6;
input 	dffe4;
input 	dffe5;
input 	pipeline_dffe_41;
input 	pipeline_dffe_31;
input 	pipeline_dffe_01;
input 	pipeline_dffe_18;
input 	pipeline_dffe_21;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[17]~q ;
wire \xordvalue[14]~q ;
wire \Add0~1_sumout ;
wire \a[16]~q ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \a[15]~q ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \a[14]~q ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \a[13]~q ;
wire \xordvalue[13]~q ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \a[12]~q ;
wire \xordvalue[12]~q ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \a[11]~q ;
wire \xordvalue[11]~q ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \a[10]~q ;
wire \xordvalue[10]~q ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \a[9]~q ;
wire \xordvalue[9]~q ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \a[8]~q ;
wire \xordvalue[8]~q ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \a[7]~q ;
wire \xordvalue[7]~q ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \a[6]~q ;
wire \xordvalue[6]~q ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \a[5]~q ;
wire \xordvalue[5]~q ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \a[4]~q ;
wire \xordvalue[4]~q ;
wire \a[0]~q ;
wire \xordvalue[0]~q ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \a[3]~q ;
wire \xordvalue[3]~q ;
wire \a[1]~q ;
wire \xordvalue[1]~q ;
wire \a[2]~q ;
wire \xordvalue[2]~q ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~65_sumout ;
wire \Add0~66 ;
wire \Add0~69_sumout ;
wire \Add0~70 ;
wire \xordvalue~0_combout ;
wire \xordvalue~1_combout ;
wire \xordvalue~2_combout ;
wire \xordvalue~3_combout ;
wire \xordvalue~4_combout ;
wire \xordvalue~5_combout ;
wire \xordvalue~6_combout ;
wire \xordvalue~7_combout ;
wire \xordvalue~8_combout ;
wire \xordvalue~9_combout ;
wire \xordvalue~10_combout ;
wire \xordvalue~11_combout ;
wire \xordvalue~12_combout ;
wire \xordvalue~13_combout ;
wire \xordvalue~14_combout ;


nco_test_lpm_add_sub_2 u0(
	.a_17(\a[17]~q ),
	.xordvalue_14(\xordvalue[14]~q ),
	.a_16(\a[16]~q ),
	.a_15(\a[15]~q ),
	.a_14(\a[14]~q ),
	.a_13(\a[13]~q ),
	.xordvalue_13(\xordvalue[13]~q ),
	.a_12(\a[12]~q ),
	.xordvalue_12(\xordvalue[12]~q ),
	.a_11(\a[11]~q ),
	.xordvalue_11(\xordvalue[11]~q ),
	.a_10(\a[10]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.a_9(\a[9]~q ),
	.xordvalue_9(\xordvalue[9]~q ),
	.a_8(\a[8]~q ),
	.xordvalue_8(\xordvalue[8]~q ),
	.a_7(\a[7]~q ),
	.xordvalue_7(\xordvalue[7]~q ),
	.a_6(\a[6]~q ),
	.xordvalue_6(\xordvalue[6]~q ),
	.a_5(\a[5]~q ),
	.xordvalue_5(\xordvalue[5]~q ),
	.a_4(\a[4]~q ),
	.xordvalue_4(\xordvalue[4]~q ),
	.a_0(\a[0]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_3(\a[3]~q ),
	.xordvalue_3(\xordvalue[3]~q ),
	.a_1(\a[1]~q ),
	.xordvalue_1(\xordvalue[1]~q ),
	.a_2(\a[2]~q ),
	.xordvalue_2(\xordvalue[2]~q ),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[17] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[17]~q ),
	.prn(vcc));
defparam \a[17] .is_wysiwyg = "true";
defparam \a[17] .power_up = "low";

dffeas \xordvalue[14] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[14]~q ),
	.prn(vcc));
defparam \xordvalue[14] .is_wysiwyg = "true";
defparam \xordvalue[14] .power_up = "low";

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_171),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h00000000000000FF;
defparam \Add0~1 .shared_arith = "off";

dffeas \a[16] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[16]~q ),
	.prn(vcc));
defparam \a[16] .is_wysiwyg = "true";
defparam \a[16] .power_up = "low";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h00000000000000FF;
defparam \Add0~5 .shared_arith = "off";

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h00000000000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h00000000000000FF;
defparam \Add0~13 .shared_arith = "off";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

dffeas \xordvalue[13] (
	.clk(clk),
	.d(\xordvalue~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[13]~q ),
	.prn(vcc));
defparam \xordvalue[13] .is_wysiwyg = "true";
defparam \xordvalue[13] .power_up = "low";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h00000000000000FF;
defparam \Add0~17 .shared_arith = "off";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

dffeas \xordvalue[12] (
	.clk(clk),
	.d(\xordvalue~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[12]~q ),
	.prn(vcc));
defparam \xordvalue[12] .is_wysiwyg = "true";
defparam \xordvalue[12] .power_up = "low";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h00000000000000FF;
defparam \Add0~21 .shared_arith = "off";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \xordvalue[11] (
	.clk(clk),
	.d(\xordvalue~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[11]~q ),
	.prn(vcc));
defparam \xordvalue[11] .is_wysiwyg = "true";
defparam \xordvalue[11] .power_up = "low";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h00000000000000FF;
defparam \Add0~25 .shared_arith = "off";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(\xordvalue~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h00000000000000FF;
defparam \Add0~29 .shared_arith = "off";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \xordvalue[9] (
	.clk(clk),
	.d(\xordvalue~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[9]~q ),
	.prn(vcc));
defparam \xordvalue[9] .is_wysiwyg = "true";
defparam \xordvalue[9] .power_up = "low";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h00000000000000FF;
defparam \Add0~33 .shared_arith = "off";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \xordvalue[8] (
	.clk(clk),
	.d(\xordvalue~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[8]~q ),
	.prn(vcc));
defparam \xordvalue[8] .is_wysiwyg = "true";
defparam \xordvalue[8] .power_up = "low";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h00000000000000FF;
defparam \Add0~37 .shared_arith = "off";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \xordvalue[7] (
	.clk(clk),
	.d(\xordvalue~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[7]~q ),
	.prn(vcc));
defparam \xordvalue[7] .is_wysiwyg = "true";
defparam \xordvalue[7] .power_up = "low";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h00000000000000FF;
defparam \Add0~41 .shared_arith = "off";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \xordvalue[6] (
	.clk(clk),
	.d(\xordvalue~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[6]~q ),
	.prn(vcc));
defparam \xordvalue[6] .is_wysiwyg = "true";
defparam \xordvalue[6] .power_up = "low";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h00000000000000FF;
defparam \Add0~45 .shared_arith = "off";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \xordvalue[5] (
	.clk(clk),
	.d(\xordvalue~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[5]~q ),
	.prn(vcc));
defparam \xordvalue[5] .is_wysiwyg = "true";
defparam \xordvalue[5] .power_up = "low";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout());
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h00000000000000FF;
defparam \Add0~49 .shared_arith = "off";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \xordvalue[4] (
	.clk(clk),
	.d(\xordvalue~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[4]~q ),
	.prn(vcc));
defparam \xordvalue[4] .is_wysiwyg = "true";
defparam \xordvalue[4] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout());
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h00000000000000FF;
defparam \Add0~53 .shared_arith = "off";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \xordvalue[3] (
	.clk(clk),
	.d(\xordvalue~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[3]~q ),
	.prn(vcc));
defparam \xordvalue[3] .is_wysiwyg = "true";
defparam \xordvalue[3] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \xordvalue[1] (
	.clk(clk),
	.d(\xordvalue~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[1]~q ),
	.prn(vcc));
defparam \xordvalue[1] .is_wysiwyg = "true";
defparam \xordvalue[1] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \xordvalue[2] (
	.clk(clk),
	.d(\xordvalue~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[2]~q ),
	.prn(vcc));
defparam \xordvalue[2] .is_wysiwyg = "true";
defparam \xordvalue[2] .power_up = "low";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe16),
	.datae(gnd),
	.dataf(!pipeline_dffe_01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout());
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~57 .shared_arith = "off";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout());
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h00000000000000FF;
defparam \Add0~61 .shared_arith = "off";

arriav_lcell_comb \Add0~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_18),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~65_sumout ),
	.cout(\Add0~66 ),
	.shareout());
defparam \Add0~65 .extended_lut = "off";
defparam \Add0~65 .lut_mask = 64'h00000000000000FF;
defparam \Add0~65 .shared_arith = "off";

arriav_lcell_comb \Add0~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~69_sumout ),
	.cout(\Add0~70 ),
	.shareout());
defparam \Add0~69 .extended_lut = "off";
defparam \Add0~69 .lut_mask = 64'h00000000000000FF;
defparam \Add0~69 .shared_arith = "off";

arriav_lcell_comb \xordvalue~0 (
	.dataa(!dffe16),
	.datab(!dffe18),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

arriav_lcell_comb \xordvalue~1 (
	.dataa(!dffe16),
	.datab(!dffe17),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~1 .extended_lut = "off";
defparam \xordvalue~1 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~1 .shared_arith = "off";

arriav_lcell_comb \xordvalue~2 (
	.dataa(!dffe16),
	.datab(!dffe161),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~2 .extended_lut = "off";
defparam \xordvalue~2 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~2 .shared_arith = "off";

arriav_lcell_comb \xordvalue~3 (
	.dataa(!dffe16),
	.datab(!dffe15),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~3 .extended_lut = "off";
defparam \xordvalue~3 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~3 .shared_arith = "off";

arriav_lcell_comb \xordvalue~4 (
	.dataa(!dffe16),
	.datab(!dffe14),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~4 .extended_lut = "off";
defparam \xordvalue~4 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~4 .shared_arith = "off";

arriav_lcell_comb \xordvalue~5 (
	.dataa(!dffe16),
	.datab(!dffe13),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~5 .extended_lut = "off";
defparam \xordvalue~5 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~5 .shared_arith = "off";

arriav_lcell_comb \xordvalue~6 (
	.dataa(!dffe16),
	.datab(!dffe12),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~6 .extended_lut = "off";
defparam \xordvalue~6 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~6 .shared_arith = "off";

arriav_lcell_comb \xordvalue~7 (
	.dataa(!dffe16),
	.datab(!dffe11),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~7 .extended_lut = "off";
defparam \xordvalue~7 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~7 .shared_arith = "off";

arriav_lcell_comb \xordvalue~8 (
	.dataa(!dffe16),
	.datab(!dffe10),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~8 .extended_lut = "off";
defparam \xordvalue~8 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~8 .shared_arith = "off";

arriav_lcell_comb \xordvalue~9 (
	.dataa(!dffe16),
	.datab(!dffe9),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~9 .extended_lut = "off";
defparam \xordvalue~9 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~9 .shared_arith = "off";

arriav_lcell_comb \xordvalue~10 (
	.dataa(!dffe16),
	.datab(!dffe8),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~10 .extended_lut = "off";
defparam \xordvalue~10 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~10 .shared_arith = "off";

arriav_lcell_comb \xordvalue~11 (
	.dataa(!dffe16),
	.datab(!dffe4),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~11 .extended_lut = "off";
defparam \xordvalue~11 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~11 .shared_arith = "off";

arriav_lcell_comb \xordvalue~12 (
	.dataa(!dffe16),
	.datab(!dffe7),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~12 .extended_lut = "off";
defparam \xordvalue~12 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~12 .shared_arith = "off";

arriav_lcell_comb \xordvalue~13 (
	.dataa(!dffe16),
	.datab(!dffe5),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~13 .extended_lut = "off";
defparam \xordvalue~13 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~13 .shared_arith = "off";

arriav_lcell_comb \xordvalue~14 (
	.dataa(!dffe16),
	.datab(!dffe6),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~14 .extended_lut = "off";
defparam \xordvalue~14 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~14 .shared_arith = "off";

endmodule

module nco_test_lpm_add_sub_2 (
	a_17,
	xordvalue_14,
	a_16,
	a_15,
	a_14,
	a_13,
	xordvalue_13,
	a_12,
	xordvalue_12,
	a_11,
	xordvalue_11,
	a_10,
	xordvalue_10,
	a_9,
	xordvalue_9,
	a_8,
	xordvalue_8,
	a_7,
	xordvalue_7,
	a_6,
	xordvalue_6,
	a_5,
	xordvalue_5,
	a_4,
	xordvalue_4,
	a_0,
	xordvalue_0,
	a_3,
	xordvalue_3,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	pipeline_dffe_17,
	pipeline_dffe_16,
	pipeline_dffe_15,
	pipeline_dffe_14,
	pipeline_dffe_13,
	pipeline_dffe_12,
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_7,
	pipeline_dffe_6,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_14;
input 	a_16;
input 	a_15;
input 	a_14;
input 	a_13;
input 	xordvalue_13;
input 	a_12;
input 	xordvalue_12;
input 	a_11;
input 	xordvalue_11;
input 	a_10;
input 	xordvalue_10;
input 	a_9;
input 	xordvalue_9;
input 	a_8;
input 	xordvalue_8;
input 	a_7;
input 	xordvalue_7;
input 	a_6;
input 	xordvalue_6;
input 	a_5;
input 	xordvalue_5;
input 	a_4;
input 	xordvalue_4;
input 	a_0;
input 	xordvalue_0;
input 	a_3;
input 	xordvalue_3;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
output 	pipeline_dffe_17;
output 	pipeline_dffe_16;
output 	pipeline_dffe_15;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_7;
output 	pipeline_dffe_6;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_add_sub_0qg auto_generated(
	.a_17(a_17),
	.xordvalue_14(xordvalue_14),
	.a_16(a_16),
	.a_15(a_15),
	.a_14(a_14),
	.a_13(a_13),
	.xordvalue_13(xordvalue_13),
	.a_12(a_12),
	.xordvalue_12(xordvalue_12),
	.a_11(a_11),
	.xordvalue_11(xordvalue_11),
	.a_10(a_10),
	.xordvalue_10(xordvalue_10),
	.a_9(a_9),
	.xordvalue_9(xordvalue_9),
	.a_8(a_8),
	.xordvalue_8(xordvalue_8),
	.a_7(a_7),
	.xordvalue_7(xordvalue_7),
	.a_6(a_6),
	.xordvalue_6(xordvalue_6),
	.a_5(a_5),
	.xordvalue_5(xordvalue_5),
	.a_4(a_4),
	.xordvalue_4(xordvalue_4),
	.a_0(a_0),
	.xordvalue_0(xordvalue_0),
	.a_3(a_3),
	.xordvalue_3(xordvalue_3),
	.a_1(a_1),
	.xordvalue_1(xordvalue_1),
	.a_2(a_2),
	.xordvalue_2(xordvalue_2),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module nco_test_add_sub_0qg (
	a_17,
	xordvalue_14,
	a_16,
	a_15,
	a_14,
	a_13,
	xordvalue_13,
	a_12,
	xordvalue_12,
	a_11,
	xordvalue_11,
	a_10,
	xordvalue_10,
	a_9,
	xordvalue_9,
	a_8,
	xordvalue_8,
	a_7,
	xordvalue_7,
	a_6,
	xordvalue_6,
	a_5,
	xordvalue_5,
	a_4,
	xordvalue_4,
	a_0,
	xordvalue_0,
	a_3,
	xordvalue_3,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	pipeline_dffe_17,
	pipeline_dffe_16,
	pipeline_dffe_15,
	pipeline_dffe_14,
	pipeline_dffe_13,
	pipeline_dffe_12,
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_7,
	pipeline_dffe_6,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_14;
input 	a_16;
input 	a_15;
input 	a_14;
input 	a_13;
input 	xordvalue_13;
input 	a_12;
input 	xordvalue_12;
input 	a_11;
input 	xordvalue_11;
input 	a_10;
input 	xordvalue_10;
input 	a_9;
input 	xordvalue_9;
input 	a_8;
input 	xordvalue_8;
input 	a_7;
input 	xordvalue_7;
input 	a_6;
input 	xordvalue_6;
input 	a_5;
input 	xordvalue_5;
input 	a_4;
input 	xordvalue_4;
input 	a_0;
input 	xordvalue_0;
input 	a_3;
input 	xordvalue_3;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
output 	pipeline_dffe_17;
output 	pipeline_dffe_16;
output 	pipeline_dffe_15;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_7;
output 	pipeline_dffe_6;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \op_1~58 ;
wire \op_1~66 ;
wire \op_1~70 ;
wire \op_1~62 ;
wire \op_1~54 ;
wire \op_1~50 ;
wire \op_1~46 ;
wire \op_1~42 ;
wire \op_1~38 ;
wire \op_1~34 ;
wire \op_1~30 ;
wire \op_1~26 ;
wire \op_1~22 ;
wire \op_1~18 ;
wire \op_1~14 ;
wire \op_1~10 ;
wire \op_1~6 ;
wire \op_1~1_sumout ;
wire \op_1~5_sumout ;
wire \op_1~9_sumout ;
wire \op_1~13_sumout ;
wire \op_1~17_sumout ;
wire \op_1~21_sumout ;
wire \op_1~25_sumout ;
wire \op_1~29_sumout ;
wire \op_1~33_sumout ;
wire \op_1~37_sumout ;
wire \op_1~41_sumout ;
wire \op_1~45_sumout ;
wire \op_1~53_sumout ;
wire \op_1~49_sumout ;
wire \op_1~57_sumout ;
wire \op_1~65_sumout ;
wire \op_1~69_sumout ;
wire \op_1~61_sumout ;


dffeas \pipeline_dffe[17] (
	.clk(clock),
	.d(\op_1~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_17),
	.prn(vcc));
defparam \pipeline_dffe[17] .is_wysiwyg = "true";
defparam \pipeline_dffe[17] .power_up = "low";

dffeas \pipeline_dffe[16] (
	.clk(clock),
	.d(\op_1~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_16),
	.prn(vcc));
defparam \pipeline_dffe[16] .is_wysiwyg = "true";
defparam \pipeline_dffe[16] .power_up = "low";

dffeas \pipeline_dffe[15] (
	.clk(clock),
	.d(\op_1~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_15),
	.prn(vcc));
defparam \pipeline_dffe[15] .is_wysiwyg = "true";
defparam \pipeline_dffe[15] .power_up = "low";

dffeas \pipeline_dffe[14] (
	.clk(clock),
	.d(\op_1~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_14),
	.prn(vcc));
defparam \pipeline_dffe[14] .is_wysiwyg = "true";
defparam \pipeline_dffe[14] .power_up = "low";

dffeas \pipeline_dffe[13] (
	.clk(clock),
	.d(\op_1~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_13),
	.prn(vcc));
defparam \pipeline_dffe[13] .is_wysiwyg = "true";
defparam \pipeline_dffe[13] .power_up = "low";

dffeas \pipeline_dffe[12] (
	.clk(clock),
	.d(\op_1~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_12),
	.prn(vcc));
defparam \pipeline_dffe[12] .is_wysiwyg = "true";
defparam \pipeline_dffe[12] .power_up = "low";

dffeas \pipeline_dffe[11] (
	.clk(clock),
	.d(\op_1~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \pipeline_dffe[11] .is_wysiwyg = "true";
defparam \pipeline_dffe[11] .power_up = "low";

dffeas \pipeline_dffe[10] (
	.clk(clock),
	.d(\op_1~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \pipeline_dffe[10] .is_wysiwyg = "true";
defparam \pipeline_dffe[10] .power_up = "low";

dffeas \pipeline_dffe[9] (
	.clk(clock),
	.d(\op_1~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \pipeline_dffe[9] .is_wysiwyg = "true";
defparam \pipeline_dffe[9] .power_up = "low";

dffeas \pipeline_dffe[8] (
	.clk(clock),
	.d(\op_1~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \pipeline_dffe[8] .is_wysiwyg = "true";
defparam \pipeline_dffe[8] .power_up = "low";

dffeas \pipeline_dffe[7] (
	.clk(clock),
	.d(\op_1~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \pipeline_dffe[7] .is_wysiwyg = "true";
defparam \pipeline_dffe[7] .power_up = "low";

dffeas \pipeline_dffe[6] (
	.clk(clock),
	.d(\op_1~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \pipeline_dffe[6] .is_wysiwyg = "true";
defparam \pipeline_dffe[6] .power_up = "low";

dffeas \pipeline_dffe[4] (
	.clk(clock),
	.d(\op_1~53_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \pipeline_dffe[4] .is_wysiwyg = "true";
defparam \pipeline_dffe[4] .power_up = "low";

dffeas \pipeline_dffe[5] (
	.clk(clock),
	.d(\op_1~49_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \pipeline_dffe[5] .is_wysiwyg = "true";
defparam \pipeline_dffe[5] .power_up = "low";

dffeas \pipeline_dffe[0] (
	.clk(clock),
	.d(\op_1~57_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_0),
	.prn(vcc));
defparam \pipeline_dffe[0] .is_wysiwyg = "true";
defparam \pipeline_dffe[0] .power_up = "low";

dffeas \pipeline_dffe[1] (
	.clk(clock),
	.d(\op_1~65_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_1),
	.prn(vcc));
defparam \pipeline_dffe[1] .is_wysiwyg = "true";
defparam \pipeline_dffe[1] .power_up = "low";

dffeas \pipeline_dffe[2] (
	.clk(clock),
	.d(\op_1~69_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \pipeline_dffe[2] .is_wysiwyg = "true";
defparam \pipeline_dffe[2] .power_up = "low";

dffeas \pipeline_dffe[3] (
	.clk(clock),
	.d(\op_1~61_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \pipeline_dffe[3] .is_wysiwyg = "true";
defparam \pipeline_dffe[3] .power_up = "low";

arriav_lcell_comb \op_1~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~57_sumout ),
	.cout(\op_1~58 ),
	.shareout());
defparam \op_1~57 .extended_lut = "off";
defparam \op_1~57 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~57 .shared_arith = "off";

arriav_lcell_comb \op_1~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_1),
	.datag(gnd),
	.cin(\op_1~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~65_sumout ),
	.cout(\op_1~66 ),
	.shareout());
defparam \op_1~65 .extended_lut = "off";
defparam \op_1~65 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~65 .shared_arith = "off";

arriav_lcell_comb \op_1~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_2),
	.datag(gnd),
	.cin(\op_1~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~69_sumout ),
	.cout(\op_1~70 ),
	.shareout());
defparam \op_1~69 .extended_lut = "off";
defparam \op_1~69 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~69 .shared_arith = "off";

arriav_lcell_comb \op_1~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_3),
	.datag(gnd),
	.cin(\op_1~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~61_sumout ),
	.cout(\op_1~62 ),
	.shareout());
defparam \op_1~61 .extended_lut = "off";
defparam \op_1~61 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~61 .shared_arith = "off";

arriav_lcell_comb \op_1~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_4),
	.datag(gnd),
	.cin(\op_1~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~53_sumout ),
	.cout(\op_1~54 ),
	.shareout());
defparam \op_1~53 .extended_lut = "off";
defparam \op_1~53 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~53 .shared_arith = "off";

arriav_lcell_comb \op_1~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_5),
	.datag(gnd),
	.cin(\op_1~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~49_sumout ),
	.cout(\op_1~50 ),
	.shareout());
defparam \op_1~49 .extended_lut = "off";
defparam \op_1~49 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~49 .shared_arith = "off";

arriav_lcell_comb \op_1~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_6),
	.datag(gnd),
	.cin(\op_1~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~45_sumout ),
	.cout(\op_1~46 ),
	.shareout());
defparam \op_1~45 .extended_lut = "off";
defparam \op_1~45 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~45 .shared_arith = "off";

arriav_lcell_comb \op_1~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_7),
	.datag(gnd),
	.cin(\op_1~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~41_sumout ),
	.cout(\op_1~42 ),
	.shareout());
defparam \op_1~41 .extended_lut = "off";
defparam \op_1~41 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~41 .shared_arith = "off";

arriav_lcell_comb \op_1~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_8),
	.datag(gnd),
	.cin(\op_1~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~37_sumout ),
	.cout(\op_1~38 ),
	.shareout());
defparam \op_1~37 .extended_lut = "off";
defparam \op_1~37 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~37 .shared_arith = "off";

arriav_lcell_comb \op_1~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_9),
	.datag(gnd),
	.cin(\op_1~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~33_sumout ),
	.cout(\op_1~34 ),
	.shareout());
defparam \op_1~33 .extended_lut = "off";
defparam \op_1~33 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~33 .shared_arith = "off";

arriav_lcell_comb \op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~29_sumout ),
	.cout(\op_1~30 ),
	.shareout());
defparam \op_1~29 .extended_lut = "off";
defparam \op_1~29 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~29 .shared_arith = "off";

arriav_lcell_comb \op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_11),
	.datag(gnd),
	.cin(\op_1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~25_sumout ),
	.cout(\op_1~26 ),
	.shareout());
defparam \op_1~25 .extended_lut = "off";
defparam \op_1~25 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~25 .shared_arith = "off";

arriav_lcell_comb \op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_12),
	.datag(gnd),
	.cin(\op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~21_sumout ),
	.cout(\op_1~22 ),
	.shareout());
defparam \op_1~21 .extended_lut = "off";
defparam \op_1~21 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~21 .shared_arith = "off";

arriav_lcell_comb \op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_13),
	.datag(gnd),
	.cin(\op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~17_sumout ),
	.cout(\op_1~18 ),
	.shareout());
defparam \op_1~17 .extended_lut = "off";
defparam \op_1~17 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~17 .shared_arith = "off";

arriav_lcell_comb \op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_14),
	.datag(gnd),
	.cin(\op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~13_sumout ),
	.cout(\op_1~14 ),
	.shareout());
defparam \op_1~13 .extended_lut = "off";
defparam \op_1~13 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~13 .shared_arith = "off";

arriav_lcell_comb \op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_14),
	.datag(gnd),
	.cin(\op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~9_sumout ),
	.cout(\op_1~10 ),
	.shareout());
defparam \op_1~9 .extended_lut = "off";
defparam \op_1~9 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~9 .shared_arith = "off";

arriav_lcell_comb \op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_16),
	.datae(gnd),
	.dataf(!xordvalue_14),
	.datag(gnd),
	.cin(\op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~5_sumout ),
	.cout(\op_1~6 ),
	.shareout());
defparam \op_1~5 .extended_lut = "off";
defparam \op_1~5 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~5 .shared_arith = "off";

arriav_lcell_comb \op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_17),
	.datae(gnd),
	.dataf(!xordvalue_14),
	.datag(gnd),
	.cin(\op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~1_sumout ),
	.cout(),
	.shareout());
defparam \op_1~1 .extended_lut = "off";
defparam \op_1~1 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~1 .shared_arith = "off";

endmodule

module nco_test_cordic_axor_1p_lpm_1 (
	sin_o_0,
	pipeline_dffe_17,
	pipeline_dffe_16,
	dffe16,
	pipeline_dffe_15,
	pipeline_dffe_171,
	dffe18,
	pipeline_dffe_14,
	pipeline_dffe_13,
	dffe17,
	pipeline_dffe_161,
	pipeline_dffe_12,
	dffe161,
	pipeline_dffe_151,
	pipeline_dffe_11,
	dffe15,
	pipeline_dffe_141,
	pipeline_dffe_10,
	dffe14,
	pipeline_dffe_131,
	pipeline_dffe_9,
	dffe13,
	pipeline_dffe_121,
	pipeline_dffe_8,
	dffe12,
	pipeline_dffe_111,
	pipeline_dffe_7,
	dffe11,
	pipeline_dffe_101,
	pipeline_dffe_6,
	dffe10,
	pipeline_dffe_5,
	pipeline_dffe_91,
	pipeline_dffe_0,
	dffe9,
	pipeline_dffe_81,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	dffe8,
	pipeline_dffe_71,
	dffe7,
	pipeline_dffe_61,
	dffe5,
	dffe6,
	pipeline_dffe_41,
	pipeline_dffe_51,
	pipeline_dffe_01,
	pipeline_dffe_18,
	pipeline_dffe_21,
	pipeline_dffe_31,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	sin_o_0;
output 	pipeline_dffe_17;
output 	pipeline_dffe_16;
input 	dffe16;
output 	pipeline_dffe_15;
input 	pipeline_dffe_171;
input 	dffe18;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
input 	dffe17;
input 	pipeline_dffe_161;
output 	pipeline_dffe_12;
input 	dffe161;
input 	pipeline_dffe_151;
output 	pipeline_dffe_11;
input 	dffe15;
input 	pipeline_dffe_141;
output 	pipeline_dffe_10;
input 	dffe14;
input 	pipeline_dffe_131;
output 	pipeline_dffe_9;
input 	dffe13;
input 	pipeline_dffe_121;
output 	pipeline_dffe_8;
input 	dffe12;
input 	pipeline_dffe_111;
output 	pipeline_dffe_7;
input 	dffe11;
input 	pipeline_dffe_101;
output 	pipeline_dffe_6;
input 	dffe10;
output 	pipeline_dffe_5;
input 	pipeline_dffe_91;
output 	pipeline_dffe_0;
input 	dffe9;
input 	pipeline_dffe_81;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
input 	dffe8;
input 	pipeline_dffe_71;
input 	dffe7;
input 	pipeline_dffe_61;
input 	dffe5;
input 	dffe6;
input 	pipeline_dffe_41;
input 	pipeline_dffe_51;
input 	pipeline_dffe_01;
input 	pipeline_dffe_18;
input 	pipeline_dffe_21;
input 	pipeline_dffe_31;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[17]~q ;
wire \xordvalue[13]~q ;
wire \Add0~1_sumout ;
wire \a[16]~q ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \a[15]~q ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \a[14]~q ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \a[13]~q ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \a[12]~q ;
wire \xordvalue[12]~q ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \a[11]~q ;
wire \xordvalue[11]~q ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \a[10]~q ;
wire \xordvalue[10]~q ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \a[9]~q ;
wire \xordvalue[9]~q ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \a[8]~q ;
wire \xordvalue[8]~q ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \a[7]~q ;
wire \xordvalue[7]~q ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \a[6]~q ;
wire \xordvalue[6]~q ;
wire \a[5]~q ;
wire \xordvalue[5]~q ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \a[0]~q ;
wire \xordvalue[0]~q ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \a[4]~q ;
wire \xordvalue[4]~q ;
wire \a[1]~q ;
wire \xordvalue[1]~q ;
wire \a[2]~q ;
wire \xordvalue[2]~q ;
wire \a[3]~q ;
wire \xordvalue[3]~q ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~65_sumout ;
wire \Add0~66 ;
wire \Add0~69_sumout ;
wire \Add0~70 ;
wire \xordvalue~0_combout ;
wire \xordvalue~1_combout ;
wire \xordvalue~2_combout ;
wire \xordvalue~3_combout ;
wire \xordvalue~4_combout ;
wire \xordvalue~5_combout ;
wire \xordvalue~6_combout ;
wire \xordvalue~7_combout ;
wire \xordvalue~8_combout ;
wire \xordvalue~9_combout ;
wire \xordvalue~10_combout ;
wire \xordvalue~11_combout ;
wire \xordvalue~12_combout ;
wire \xordvalue~13_combout ;


nco_test_lpm_add_sub_3 u0(
	.a_17(\a[17]~q ),
	.xordvalue_13(\xordvalue[13]~q ),
	.a_16(\a[16]~q ),
	.a_15(\a[15]~q ),
	.a_14(\a[14]~q ),
	.a_13(\a[13]~q ),
	.a_12(\a[12]~q ),
	.xordvalue_12(\xordvalue[12]~q ),
	.a_11(\a[11]~q ),
	.xordvalue_11(\xordvalue[11]~q ),
	.a_10(\a[10]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.a_9(\a[9]~q ),
	.xordvalue_9(\xordvalue[9]~q ),
	.a_8(\a[8]~q ),
	.xordvalue_8(\xordvalue[8]~q ),
	.a_7(\a[7]~q ),
	.xordvalue_7(\xordvalue[7]~q ),
	.a_6(\a[6]~q ),
	.xordvalue_6(\xordvalue[6]~q ),
	.a_5(\a[5]~q ),
	.xordvalue_5(\xordvalue[5]~q ),
	.a_0(\a[0]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_4(\a[4]~q ),
	.xordvalue_4(\xordvalue[4]~q ),
	.a_1(\a[1]~q ),
	.xordvalue_1(\xordvalue[1]~q ),
	.a_2(\a[2]~q ),
	.xordvalue_2(\xordvalue[2]~q ),
	.a_3(\a[3]~q ),
	.xordvalue_3(\xordvalue[3]~q ),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[17] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[17]~q ),
	.prn(vcc));
defparam \a[17] .is_wysiwyg = "true";
defparam \a[17] .power_up = "low";

dffeas \xordvalue[13] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[13]~q ),
	.prn(vcc));
defparam \xordvalue[13] .is_wysiwyg = "true";
defparam \xordvalue[13] .power_up = "low";

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_171),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h00000000000000FF;
defparam \Add0~1 .shared_arith = "off";

dffeas \a[16] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[16]~q ),
	.prn(vcc));
defparam \a[16] .is_wysiwyg = "true";
defparam \a[16] .power_up = "low";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h00000000000000FF;
defparam \Add0~5 .shared_arith = "off";

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h00000000000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h00000000000000FF;
defparam \Add0~13 .shared_arith = "off";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h00000000000000FF;
defparam \Add0~17 .shared_arith = "off";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

dffeas \xordvalue[12] (
	.clk(clk),
	.d(\xordvalue~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[12]~q ),
	.prn(vcc));
defparam \xordvalue[12] .is_wysiwyg = "true";
defparam \xordvalue[12] .power_up = "low";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h00000000000000FF;
defparam \Add0~21 .shared_arith = "off";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \xordvalue[11] (
	.clk(clk),
	.d(\xordvalue~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[11]~q ),
	.prn(vcc));
defparam \xordvalue[11] .is_wysiwyg = "true";
defparam \xordvalue[11] .power_up = "low";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h00000000000000FF;
defparam \Add0~25 .shared_arith = "off";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(\xordvalue~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h00000000000000FF;
defparam \Add0~29 .shared_arith = "off";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \xordvalue[9] (
	.clk(clk),
	.d(\xordvalue~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[9]~q ),
	.prn(vcc));
defparam \xordvalue[9] .is_wysiwyg = "true";
defparam \xordvalue[9] .power_up = "low";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h00000000000000FF;
defparam \Add0~33 .shared_arith = "off";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \xordvalue[8] (
	.clk(clk),
	.d(\xordvalue~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[8]~q ),
	.prn(vcc));
defparam \xordvalue[8] .is_wysiwyg = "true";
defparam \xordvalue[8] .power_up = "low";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h00000000000000FF;
defparam \Add0~37 .shared_arith = "off";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \xordvalue[7] (
	.clk(clk),
	.d(\xordvalue~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[7]~q ),
	.prn(vcc));
defparam \xordvalue[7] .is_wysiwyg = "true";
defparam \xordvalue[7] .power_up = "low";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h00000000000000FF;
defparam \Add0~41 .shared_arith = "off";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \xordvalue[6] (
	.clk(clk),
	.d(\xordvalue~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[6]~q ),
	.prn(vcc));
defparam \xordvalue[6] .is_wysiwyg = "true";
defparam \xordvalue[6] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \xordvalue[5] (
	.clk(clk),
	.d(\xordvalue~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[5]~q ),
	.prn(vcc));
defparam \xordvalue[5] .is_wysiwyg = "true";
defparam \xordvalue[5] .power_up = "low";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h00000000000000FF;
defparam \Add0~45 .shared_arith = "off";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout());
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h00000000000000FF;
defparam \Add0~49 .shared_arith = "off";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \xordvalue[4] (
	.clk(clk),
	.d(\xordvalue~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[4]~q ),
	.prn(vcc));
defparam \xordvalue[4] .is_wysiwyg = "true";
defparam \xordvalue[4] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \xordvalue[1] (
	.clk(clk),
	.d(\xordvalue~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[1]~q ),
	.prn(vcc));
defparam \xordvalue[1] .is_wysiwyg = "true";
defparam \xordvalue[1] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \xordvalue[2] (
	.clk(clk),
	.d(\xordvalue~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[2]~q ),
	.prn(vcc));
defparam \xordvalue[2] .is_wysiwyg = "true";
defparam \xordvalue[2] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \xordvalue[3] (
	.clk(clk),
	.d(\xordvalue~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[3]~q ),
	.prn(vcc));
defparam \xordvalue[3] .is_wysiwyg = "true";
defparam \xordvalue[3] .power_up = "low";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe16),
	.datae(gnd),
	.dataf(!pipeline_dffe_01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout());
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~53 .shared_arith = "off";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout());
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h00000000000000FF;
defparam \Add0~57 .shared_arith = "off";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_18),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout());
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h00000000000000FF;
defparam \Add0~61 .shared_arith = "off";

arriav_lcell_comb \Add0~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~65_sumout ),
	.cout(\Add0~66 ),
	.shareout());
defparam \Add0~65 .extended_lut = "off";
defparam \Add0~65 .lut_mask = 64'h00000000000000FF;
defparam \Add0~65 .shared_arith = "off";

arriav_lcell_comb \Add0~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~69_sumout ),
	.cout(\Add0~70 ),
	.shareout());
defparam \Add0~69 .extended_lut = "off";
defparam \Add0~69 .lut_mask = 64'h00000000000000FF;
defparam \Add0~69 .shared_arith = "off";

arriav_lcell_comb \xordvalue~0 (
	.dataa(!dffe18),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

arriav_lcell_comb \xordvalue~1 (
	.dataa(!dffe17),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~1 .extended_lut = "off";
defparam \xordvalue~1 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~1 .shared_arith = "off";

arriav_lcell_comb \xordvalue~2 (
	.dataa(!dffe161),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~2 .extended_lut = "off";
defparam \xordvalue~2 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~2 .shared_arith = "off";

arriav_lcell_comb \xordvalue~3 (
	.dataa(!dffe15),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~3 .extended_lut = "off";
defparam \xordvalue~3 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~3 .shared_arith = "off";

arriav_lcell_comb \xordvalue~4 (
	.dataa(!dffe14),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~4 .extended_lut = "off";
defparam \xordvalue~4 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~4 .shared_arith = "off";

arriav_lcell_comb \xordvalue~5 (
	.dataa(!dffe13),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~5 .extended_lut = "off";
defparam \xordvalue~5 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~5 .shared_arith = "off";

arriav_lcell_comb \xordvalue~6 (
	.dataa(!dffe12),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~6 .extended_lut = "off";
defparam \xordvalue~6 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~6 .shared_arith = "off";

arriav_lcell_comb \xordvalue~7 (
	.dataa(!dffe11),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~7 .extended_lut = "off";
defparam \xordvalue~7 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~7 .shared_arith = "off";

arriav_lcell_comb \xordvalue~8 (
	.dataa(!dffe10),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~8 .extended_lut = "off";
defparam \xordvalue~8 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~8 .shared_arith = "off";

arriav_lcell_comb \xordvalue~9 (
	.dataa(!dffe5),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~9 .extended_lut = "off";
defparam \xordvalue~9 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~9 .shared_arith = "off";

arriav_lcell_comb \xordvalue~10 (
	.dataa(!dffe9),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~10 .extended_lut = "off";
defparam \xordvalue~10 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~10 .shared_arith = "off";

arriav_lcell_comb \xordvalue~11 (
	.dataa(!dffe6),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~11 .extended_lut = "off";
defparam \xordvalue~11 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~11 .shared_arith = "off";

arriav_lcell_comb \xordvalue~12 (
	.dataa(!dffe7),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~12 .extended_lut = "off";
defparam \xordvalue~12 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~12 .shared_arith = "off";

arriav_lcell_comb \xordvalue~13 (
	.dataa(!dffe8),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~13 .extended_lut = "off";
defparam \xordvalue~13 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~13 .shared_arith = "off";

endmodule

module nco_test_lpm_add_sub_3 (
	a_17,
	xordvalue_13,
	a_16,
	a_15,
	a_14,
	a_13,
	a_12,
	xordvalue_12,
	a_11,
	xordvalue_11,
	a_10,
	xordvalue_10,
	a_9,
	xordvalue_9,
	a_8,
	xordvalue_8,
	a_7,
	xordvalue_7,
	a_6,
	xordvalue_6,
	a_5,
	xordvalue_5,
	a_0,
	xordvalue_0,
	a_4,
	xordvalue_4,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	pipeline_dffe_17,
	pipeline_dffe_16,
	pipeline_dffe_15,
	pipeline_dffe_14,
	pipeline_dffe_13,
	pipeline_dffe_12,
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_7,
	pipeline_dffe_6,
	pipeline_dffe_5,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_13;
input 	a_16;
input 	a_15;
input 	a_14;
input 	a_13;
input 	a_12;
input 	xordvalue_12;
input 	a_11;
input 	xordvalue_11;
input 	a_10;
input 	xordvalue_10;
input 	a_9;
input 	xordvalue_9;
input 	a_8;
input 	xordvalue_8;
input 	a_7;
input 	xordvalue_7;
input 	a_6;
input 	xordvalue_6;
input 	a_5;
input 	xordvalue_5;
input 	a_0;
input 	xordvalue_0;
input 	a_4;
input 	xordvalue_4;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
output 	pipeline_dffe_17;
output 	pipeline_dffe_16;
output 	pipeline_dffe_15;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_7;
output 	pipeline_dffe_6;
output 	pipeline_dffe_5;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_add_sub_0qg_1 auto_generated(
	.a_17(a_17),
	.xordvalue_13(xordvalue_13),
	.a_16(a_16),
	.a_15(a_15),
	.a_14(a_14),
	.a_13(a_13),
	.a_12(a_12),
	.xordvalue_12(xordvalue_12),
	.a_11(a_11),
	.xordvalue_11(xordvalue_11),
	.a_10(a_10),
	.xordvalue_10(xordvalue_10),
	.a_9(a_9),
	.xordvalue_9(xordvalue_9),
	.a_8(a_8),
	.xordvalue_8(xordvalue_8),
	.a_7(a_7),
	.xordvalue_7(xordvalue_7),
	.a_6(a_6),
	.xordvalue_6(xordvalue_6),
	.a_5(a_5),
	.xordvalue_5(xordvalue_5),
	.a_0(a_0),
	.xordvalue_0(xordvalue_0),
	.a_4(a_4),
	.xordvalue_4(xordvalue_4),
	.a_1(a_1),
	.xordvalue_1(xordvalue_1),
	.a_2(a_2),
	.xordvalue_2(xordvalue_2),
	.a_3(a_3),
	.xordvalue_3(xordvalue_3),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module nco_test_add_sub_0qg_1 (
	a_17,
	xordvalue_13,
	a_16,
	a_15,
	a_14,
	a_13,
	a_12,
	xordvalue_12,
	a_11,
	xordvalue_11,
	a_10,
	xordvalue_10,
	a_9,
	xordvalue_9,
	a_8,
	xordvalue_8,
	a_7,
	xordvalue_7,
	a_6,
	xordvalue_6,
	a_5,
	xordvalue_5,
	a_0,
	xordvalue_0,
	a_4,
	xordvalue_4,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	pipeline_dffe_17,
	pipeline_dffe_16,
	pipeline_dffe_15,
	pipeline_dffe_14,
	pipeline_dffe_13,
	pipeline_dffe_12,
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_7,
	pipeline_dffe_6,
	pipeline_dffe_5,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_13;
input 	a_16;
input 	a_15;
input 	a_14;
input 	a_13;
input 	a_12;
input 	xordvalue_12;
input 	a_11;
input 	xordvalue_11;
input 	a_10;
input 	xordvalue_10;
input 	a_9;
input 	xordvalue_9;
input 	a_8;
input 	xordvalue_8;
input 	a_7;
input 	xordvalue_7;
input 	a_6;
input 	xordvalue_6;
input 	a_5;
input 	xordvalue_5;
input 	a_0;
input 	xordvalue_0;
input 	a_4;
input 	xordvalue_4;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
output 	pipeline_dffe_17;
output 	pipeline_dffe_16;
output 	pipeline_dffe_15;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_7;
output 	pipeline_dffe_6;
output 	pipeline_dffe_5;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \op_1~54 ;
wire \op_1~62 ;
wire \op_1~66 ;
wire \op_1~70 ;
wire \op_1~58 ;
wire \op_1~50 ;
wire \op_1~46 ;
wire \op_1~42 ;
wire \op_1~38 ;
wire \op_1~34 ;
wire \op_1~30 ;
wire \op_1~26 ;
wire \op_1~22 ;
wire \op_1~18 ;
wire \op_1~14 ;
wire \op_1~10 ;
wire \op_1~6 ;
wire \op_1~1_sumout ;
wire \op_1~5_sumout ;
wire \op_1~9_sumout ;
wire \op_1~13_sumout ;
wire \op_1~17_sumout ;
wire \op_1~21_sumout ;
wire \op_1~25_sumout ;
wire \op_1~29_sumout ;
wire \op_1~33_sumout ;
wire \op_1~37_sumout ;
wire \op_1~41_sumout ;
wire \op_1~45_sumout ;
wire \op_1~49_sumout ;
wire \op_1~53_sumout ;
wire \op_1~61_sumout ;
wire \op_1~65_sumout ;
wire \op_1~69_sumout ;
wire \op_1~57_sumout ;


dffeas \pipeline_dffe[17] (
	.clk(clock),
	.d(\op_1~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_17),
	.prn(vcc));
defparam \pipeline_dffe[17] .is_wysiwyg = "true";
defparam \pipeline_dffe[17] .power_up = "low";

dffeas \pipeline_dffe[16] (
	.clk(clock),
	.d(\op_1~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_16),
	.prn(vcc));
defparam \pipeline_dffe[16] .is_wysiwyg = "true";
defparam \pipeline_dffe[16] .power_up = "low";

dffeas \pipeline_dffe[15] (
	.clk(clock),
	.d(\op_1~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_15),
	.prn(vcc));
defparam \pipeline_dffe[15] .is_wysiwyg = "true";
defparam \pipeline_dffe[15] .power_up = "low";

dffeas \pipeline_dffe[14] (
	.clk(clock),
	.d(\op_1~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_14),
	.prn(vcc));
defparam \pipeline_dffe[14] .is_wysiwyg = "true";
defparam \pipeline_dffe[14] .power_up = "low";

dffeas \pipeline_dffe[13] (
	.clk(clock),
	.d(\op_1~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_13),
	.prn(vcc));
defparam \pipeline_dffe[13] .is_wysiwyg = "true";
defparam \pipeline_dffe[13] .power_up = "low";

dffeas \pipeline_dffe[12] (
	.clk(clock),
	.d(\op_1~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_12),
	.prn(vcc));
defparam \pipeline_dffe[12] .is_wysiwyg = "true";
defparam \pipeline_dffe[12] .power_up = "low";

dffeas \pipeline_dffe[11] (
	.clk(clock),
	.d(\op_1~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \pipeline_dffe[11] .is_wysiwyg = "true";
defparam \pipeline_dffe[11] .power_up = "low";

dffeas \pipeline_dffe[10] (
	.clk(clock),
	.d(\op_1~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \pipeline_dffe[10] .is_wysiwyg = "true";
defparam \pipeline_dffe[10] .power_up = "low";

dffeas \pipeline_dffe[9] (
	.clk(clock),
	.d(\op_1~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \pipeline_dffe[9] .is_wysiwyg = "true";
defparam \pipeline_dffe[9] .power_up = "low";

dffeas \pipeline_dffe[8] (
	.clk(clock),
	.d(\op_1~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \pipeline_dffe[8] .is_wysiwyg = "true";
defparam \pipeline_dffe[8] .power_up = "low";

dffeas \pipeline_dffe[7] (
	.clk(clock),
	.d(\op_1~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \pipeline_dffe[7] .is_wysiwyg = "true";
defparam \pipeline_dffe[7] .power_up = "low";

dffeas \pipeline_dffe[6] (
	.clk(clock),
	.d(\op_1~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \pipeline_dffe[6] .is_wysiwyg = "true";
defparam \pipeline_dffe[6] .power_up = "low";

dffeas \pipeline_dffe[5] (
	.clk(clock),
	.d(\op_1~49_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \pipeline_dffe[5] .is_wysiwyg = "true";
defparam \pipeline_dffe[5] .power_up = "low";

dffeas \pipeline_dffe[0] (
	.clk(clock),
	.d(\op_1~53_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_0),
	.prn(vcc));
defparam \pipeline_dffe[0] .is_wysiwyg = "true";
defparam \pipeline_dffe[0] .power_up = "low";

dffeas \pipeline_dffe[1] (
	.clk(clock),
	.d(\op_1~61_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_1),
	.prn(vcc));
defparam \pipeline_dffe[1] .is_wysiwyg = "true";
defparam \pipeline_dffe[1] .power_up = "low";

dffeas \pipeline_dffe[2] (
	.clk(clock),
	.d(\op_1~65_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \pipeline_dffe[2] .is_wysiwyg = "true";
defparam \pipeline_dffe[2] .power_up = "low";

dffeas \pipeline_dffe[3] (
	.clk(clock),
	.d(\op_1~69_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \pipeline_dffe[3] .is_wysiwyg = "true";
defparam \pipeline_dffe[3] .power_up = "low";

dffeas \pipeline_dffe[4] (
	.clk(clock),
	.d(\op_1~57_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \pipeline_dffe[4] .is_wysiwyg = "true";
defparam \pipeline_dffe[4] .power_up = "low";

arriav_lcell_comb \op_1~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~53_sumout ),
	.cout(\op_1~54 ),
	.shareout());
defparam \op_1~53 .extended_lut = "off";
defparam \op_1~53 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~53 .shared_arith = "off";

arriav_lcell_comb \op_1~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_1),
	.datag(gnd),
	.cin(\op_1~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~61_sumout ),
	.cout(\op_1~62 ),
	.shareout());
defparam \op_1~61 .extended_lut = "off";
defparam \op_1~61 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~61 .shared_arith = "off";

arriav_lcell_comb \op_1~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_2),
	.datag(gnd),
	.cin(\op_1~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~65_sumout ),
	.cout(\op_1~66 ),
	.shareout());
defparam \op_1~65 .extended_lut = "off";
defparam \op_1~65 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~65 .shared_arith = "off";

arriav_lcell_comb \op_1~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_3),
	.datag(gnd),
	.cin(\op_1~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~69_sumout ),
	.cout(\op_1~70 ),
	.shareout());
defparam \op_1~69 .extended_lut = "off";
defparam \op_1~69 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~69 .shared_arith = "off";

arriav_lcell_comb \op_1~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_4),
	.datag(gnd),
	.cin(\op_1~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~57_sumout ),
	.cout(\op_1~58 ),
	.shareout());
defparam \op_1~57 .extended_lut = "off";
defparam \op_1~57 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~57 .shared_arith = "off";

arriav_lcell_comb \op_1~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_5),
	.datag(gnd),
	.cin(\op_1~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~49_sumout ),
	.cout(\op_1~50 ),
	.shareout());
defparam \op_1~49 .extended_lut = "off";
defparam \op_1~49 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~49 .shared_arith = "off";

arriav_lcell_comb \op_1~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_6),
	.datag(gnd),
	.cin(\op_1~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~45_sumout ),
	.cout(\op_1~46 ),
	.shareout());
defparam \op_1~45 .extended_lut = "off";
defparam \op_1~45 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~45 .shared_arith = "off";

arriav_lcell_comb \op_1~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_7),
	.datag(gnd),
	.cin(\op_1~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~41_sumout ),
	.cout(\op_1~42 ),
	.shareout());
defparam \op_1~41 .extended_lut = "off";
defparam \op_1~41 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~41 .shared_arith = "off";

arriav_lcell_comb \op_1~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_8),
	.datag(gnd),
	.cin(\op_1~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~37_sumout ),
	.cout(\op_1~38 ),
	.shareout());
defparam \op_1~37 .extended_lut = "off";
defparam \op_1~37 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~37 .shared_arith = "off";

arriav_lcell_comb \op_1~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_9),
	.datag(gnd),
	.cin(\op_1~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~33_sumout ),
	.cout(\op_1~34 ),
	.shareout());
defparam \op_1~33 .extended_lut = "off";
defparam \op_1~33 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~33 .shared_arith = "off";

arriav_lcell_comb \op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~29_sumout ),
	.cout(\op_1~30 ),
	.shareout());
defparam \op_1~29 .extended_lut = "off";
defparam \op_1~29 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~29 .shared_arith = "off";

arriav_lcell_comb \op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_11),
	.datag(gnd),
	.cin(\op_1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~25_sumout ),
	.cout(\op_1~26 ),
	.shareout());
defparam \op_1~25 .extended_lut = "off";
defparam \op_1~25 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~25 .shared_arith = "off";

arriav_lcell_comb \op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_12),
	.datag(gnd),
	.cin(\op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~21_sumout ),
	.cout(\op_1~22 ),
	.shareout());
defparam \op_1~21 .extended_lut = "off";
defparam \op_1~21 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~21 .shared_arith = "off";

arriav_lcell_comb \op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_13),
	.datag(gnd),
	.cin(\op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~17_sumout ),
	.cout(\op_1~18 ),
	.shareout());
defparam \op_1~17 .extended_lut = "off";
defparam \op_1~17 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~17 .shared_arith = "off";

arriav_lcell_comb \op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_13),
	.datag(gnd),
	.cin(\op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~13_sumout ),
	.cout(\op_1~14 ),
	.shareout());
defparam \op_1~13 .extended_lut = "off";
defparam \op_1~13 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~13 .shared_arith = "off";

arriav_lcell_comb \op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_13),
	.datag(gnd),
	.cin(\op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~9_sumout ),
	.cout(\op_1~10 ),
	.shareout());
defparam \op_1~9 .extended_lut = "off";
defparam \op_1~9 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~9 .shared_arith = "off";

arriav_lcell_comb \op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_16),
	.datae(gnd),
	.dataf(!xordvalue_13),
	.datag(gnd),
	.cin(\op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~5_sumout ),
	.cout(\op_1~6 ),
	.shareout());
defparam \op_1~5 .extended_lut = "off";
defparam \op_1~5 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~5 .shared_arith = "off";

arriav_lcell_comb \op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_17),
	.datae(gnd),
	.dataf(!xordvalue_13),
	.datag(gnd),
	.cin(\op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~1_sumout ),
	.cout(),
	.shareout());
defparam \op_1~1 .extended_lut = "off";
defparam \op_1~1 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~1 .shared_arith = "off";

endmodule

module nco_test_cordic_axor_1p_lpm_2 (
	sin_o_0,
	pipeline_dffe_17,
	pipeline_dffe_16,
	dffe16,
	dffe18,
	pipeline_dffe_15,
	pipeline_dffe_171,
	pipeline_dffe_14,
	pipeline_dffe_161,
	pipeline_dffe_13,
	dffe17,
	pipeline_dffe_151,
	pipeline_dffe_12,
	dffe161,
	pipeline_dffe_141,
	pipeline_dffe_11,
	dffe15,
	pipeline_dffe_131,
	pipeline_dffe_10,
	dffe14,
	pipeline_dffe_121,
	pipeline_dffe_9,
	dffe13,
	pipeline_dffe_111,
	pipeline_dffe_8,
	dffe12,
	pipeline_dffe_101,
	pipeline_dffe_6,
	pipeline_dffe_7,
	dffe11,
	pipeline_dffe_0,
	pipeline_dffe_91,
	dffe10,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_81,
	dffe9,
	pipeline_dffe_71,
	dffe8,
	dffe6,
	dffe7,
	pipeline_dffe_61,
	pipeline_dffe_51,
	pipeline_dffe_01,
	pipeline_dffe_18,
	pipeline_dffe_21,
	pipeline_dffe_31,
	pipeline_dffe_41,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	sin_o_0;
output 	pipeline_dffe_17;
output 	pipeline_dffe_16;
input 	dffe16;
input 	dffe18;
output 	pipeline_dffe_15;
input 	pipeline_dffe_171;
output 	pipeline_dffe_14;
input 	pipeline_dffe_161;
output 	pipeline_dffe_13;
input 	dffe17;
input 	pipeline_dffe_151;
output 	pipeline_dffe_12;
input 	dffe161;
input 	pipeline_dffe_141;
output 	pipeline_dffe_11;
input 	dffe15;
input 	pipeline_dffe_131;
output 	pipeline_dffe_10;
input 	dffe14;
input 	pipeline_dffe_121;
output 	pipeline_dffe_9;
input 	dffe13;
input 	pipeline_dffe_111;
output 	pipeline_dffe_8;
input 	dffe12;
input 	pipeline_dffe_101;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
input 	dffe11;
output 	pipeline_dffe_0;
input 	pipeline_dffe_91;
input 	dffe10;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
input 	pipeline_dffe_81;
input 	dffe9;
input 	pipeline_dffe_71;
input 	dffe8;
input 	dffe6;
input 	dffe7;
input 	pipeline_dffe_61;
input 	pipeline_dffe_51;
input 	pipeline_dffe_01;
input 	pipeline_dffe_18;
input 	pipeline_dffe_21;
input 	pipeline_dffe_31;
input 	pipeline_dffe_41;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[17]~q ;
wire \xordvalue[12]~q ;
wire \Add0~1_sumout ;
wire \a[16]~q ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \a[15]~q ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \a[14]~q ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \a[13]~q ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \a[12]~q ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \a[11]~q ;
wire \xordvalue[11]~q ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \a[10]~q ;
wire \xordvalue[10]~q ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \a[9]~q ;
wire \xordvalue[9]~q ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \a[8]~q ;
wire \xordvalue[8]~q ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \a[7]~q ;
wire \xordvalue[7]~q ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \a[6]~q ;
wire \xordvalue[6]~q ;
wire \a[0]~q ;
wire \xordvalue[0]~q ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \a[5]~q ;
wire \xordvalue[5]~q ;
wire \a[1]~q ;
wire \xordvalue[1]~q ;
wire \a[2]~q ;
wire \xordvalue[2]~q ;
wire \a[3]~q ;
wire \xordvalue[3]~q ;
wire \a[4]~q ;
wire \xordvalue[4]~q ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~65_sumout ;
wire \Add0~66 ;
wire \Add0~69_sumout ;
wire \Add0~70 ;
wire \xordvalue~0_combout ;
wire \xordvalue~1_combout ;
wire \xordvalue~2_combout ;
wire \xordvalue~3_combout ;
wire \xordvalue~4_combout ;
wire \xordvalue~5_combout ;
wire \xordvalue~6_combout ;
wire \xordvalue~7_combout ;
wire \xordvalue~8_combout ;
wire \xordvalue~9_combout ;
wire \xordvalue~10_combout ;
wire \xordvalue~11_combout ;
wire \xordvalue~12_combout ;


nco_test_lpm_add_sub_4 u0(
	.a_17(\a[17]~q ),
	.xordvalue_12(\xordvalue[12]~q ),
	.a_16(\a[16]~q ),
	.a_15(\a[15]~q ),
	.a_14(\a[14]~q ),
	.a_13(\a[13]~q ),
	.a_12(\a[12]~q ),
	.a_11(\a[11]~q ),
	.xordvalue_11(\xordvalue[11]~q ),
	.a_10(\a[10]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.a_9(\a[9]~q ),
	.xordvalue_9(\xordvalue[9]~q ),
	.a_8(\a[8]~q ),
	.xordvalue_8(\xordvalue[8]~q ),
	.a_7(\a[7]~q ),
	.xordvalue_7(\xordvalue[7]~q ),
	.a_6(\a[6]~q ),
	.xordvalue_6(\xordvalue[6]~q ),
	.a_0(\a[0]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_5(\a[5]~q ),
	.xordvalue_5(\xordvalue[5]~q ),
	.a_1(\a[1]~q ),
	.xordvalue_1(\xordvalue[1]~q ),
	.a_2(\a[2]~q ),
	.xordvalue_2(\xordvalue[2]~q ),
	.a_3(\a[3]~q ),
	.xordvalue_3(\xordvalue[3]~q ),
	.a_4(\a[4]~q ),
	.xordvalue_4(\xordvalue[4]~q ),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[17] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[17]~q ),
	.prn(vcc));
defparam \a[17] .is_wysiwyg = "true";
defparam \a[17] .power_up = "low";

dffeas \xordvalue[12] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[12]~q ),
	.prn(vcc));
defparam \xordvalue[12] .is_wysiwyg = "true";
defparam \xordvalue[12] .power_up = "low";

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_171),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h00000000000000FF;
defparam \Add0~1 .shared_arith = "off";

dffeas \a[16] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[16]~q ),
	.prn(vcc));
defparam \a[16] .is_wysiwyg = "true";
defparam \a[16] .power_up = "low";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h00000000000000FF;
defparam \Add0~5 .shared_arith = "off";

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h00000000000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h00000000000000FF;
defparam \Add0~13 .shared_arith = "off";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h00000000000000FF;
defparam \Add0~17 .shared_arith = "off";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h00000000000000FF;
defparam \Add0~21 .shared_arith = "off";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \xordvalue[11] (
	.clk(clk),
	.d(\xordvalue~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[11]~q ),
	.prn(vcc));
defparam \xordvalue[11] .is_wysiwyg = "true";
defparam \xordvalue[11] .power_up = "low";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h00000000000000FF;
defparam \Add0~25 .shared_arith = "off";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(\xordvalue~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h00000000000000FF;
defparam \Add0~29 .shared_arith = "off";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \xordvalue[9] (
	.clk(clk),
	.d(\xordvalue~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[9]~q ),
	.prn(vcc));
defparam \xordvalue[9] .is_wysiwyg = "true";
defparam \xordvalue[9] .power_up = "low";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h00000000000000FF;
defparam \Add0~33 .shared_arith = "off";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \xordvalue[8] (
	.clk(clk),
	.d(\xordvalue~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[8]~q ),
	.prn(vcc));
defparam \xordvalue[8] .is_wysiwyg = "true";
defparam \xordvalue[8] .power_up = "low";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h00000000000000FF;
defparam \Add0~37 .shared_arith = "off";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \xordvalue[7] (
	.clk(clk),
	.d(\xordvalue~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[7]~q ),
	.prn(vcc));
defparam \xordvalue[7] .is_wysiwyg = "true";
defparam \xordvalue[7] .power_up = "low";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h00000000000000FF;
defparam \Add0~41 .shared_arith = "off";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \xordvalue[6] (
	.clk(clk),
	.d(\xordvalue~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[6]~q ),
	.prn(vcc));
defparam \xordvalue[6] .is_wysiwyg = "true";
defparam \xordvalue[6] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h00000000000000FF;
defparam \Add0~45 .shared_arith = "off";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \xordvalue[5] (
	.clk(clk),
	.d(\xordvalue~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[5]~q ),
	.prn(vcc));
defparam \xordvalue[5] .is_wysiwyg = "true";
defparam \xordvalue[5] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \xordvalue[1] (
	.clk(clk),
	.d(\xordvalue~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[1]~q ),
	.prn(vcc));
defparam \xordvalue[1] .is_wysiwyg = "true";
defparam \xordvalue[1] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \xordvalue[2] (
	.clk(clk),
	.d(\xordvalue~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[2]~q ),
	.prn(vcc));
defparam \xordvalue[2] .is_wysiwyg = "true";
defparam \xordvalue[2] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \xordvalue[3] (
	.clk(clk),
	.d(\xordvalue~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[3]~q ),
	.prn(vcc));
defparam \xordvalue[3] .is_wysiwyg = "true";
defparam \xordvalue[3] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \xordvalue[4] (
	.clk(clk),
	.d(\xordvalue~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[4]~q ),
	.prn(vcc));
defparam \xordvalue[4] .is_wysiwyg = "true";
defparam \xordvalue[4] .power_up = "low";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe16),
	.datae(gnd),
	.dataf(!pipeline_dffe_01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout());
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~49 .shared_arith = "off";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout());
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h00000000000000FF;
defparam \Add0~53 .shared_arith = "off";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_18),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout());
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h00000000000000FF;
defparam \Add0~57 .shared_arith = "off";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout());
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h00000000000000FF;
defparam \Add0~61 .shared_arith = "off";

arriav_lcell_comb \Add0~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~65_sumout ),
	.cout(\Add0~66 ),
	.shareout());
defparam \Add0~65 .extended_lut = "off";
defparam \Add0~65 .lut_mask = 64'h00000000000000FF;
defparam \Add0~65 .shared_arith = "off";

arriav_lcell_comb \Add0~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~69_sumout ),
	.cout(\Add0~70 ),
	.shareout());
defparam \Add0~69 .extended_lut = "off";
defparam \Add0~69 .lut_mask = 64'h00000000000000FF;
defparam \Add0~69 .shared_arith = "off";

arriav_lcell_comb \xordvalue~0 (
	.dataa(!dffe16),
	.datab(!dffe18),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

arriav_lcell_comb \xordvalue~1 (
	.dataa(!dffe16),
	.datab(!dffe17),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~1 .extended_lut = "off";
defparam \xordvalue~1 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~1 .shared_arith = "off";

arriav_lcell_comb \xordvalue~2 (
	.dataa(!dffe16),
	.datab(!dffe161),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~2 .extended_lut = "off";
defparam \xordvalue~2 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~2 .shared_arith = "off";

arriav_lcell_comb \xordvalue~3 (
	.dataa(!dffe16),
	.datab(!dffe15),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~3 .extended_lut = "off";
defparam \xordvalue~3 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~3 .shared_arith = "off";

arriav_lcell_comb \xordvalue~4 (
	.dataa(!dffe16),
	.datab(!dffe14),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~4 .extended_lut = "off";
defparam \xordvalue~4 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~4 .shared_arith = "off";

arriav_lcell_comb \xordvalue~5 (
	.dataa(!dffe16),
	.datab(!dffe13),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~5 .extended_lut = "off";
defparam \xordvalue~5 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~5 .shared_arith = "off";

arriav_lcell_comb \xordvalue~6 (
	.dataa(!dffe16),
	.datab(!dffe12),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~6 .extended_lut = "off";
defparam \xordvalue~6 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~6 .shared_arith = "off";

arriav_lcell_comb \xordvalue~7 (
	.dataa(!dffe16),
	.datab(!dffe6),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~7 .extended_lut = "off";
defparam \xordvalue~7 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~7 .shared_arith = "off";

arriav_lcell_comb \xordvalue~8 (
	.dataa(!dffe16),
	.datab(!dffe11),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~8 .extended_lut = "off";
defparam \xordvalue~8 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~8 .shared_arith = "off";

arriav_lcell_comb \xordvalue~9 (
	.dataa(!dffe16),
	.datab(!dffe7),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~9 .extended_lut = "off";
defparam \xordvalue~9 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~9 .shared_arith = "off";

arriav_lcell_comb \xordvalue~10 (
	.dataa(!dffe16),
	.datab(!dffe8),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~10 .extended_lut = "off";
defparam \xordvalue~10 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~10 .shared_arith = "off";

arriav_lcell_comb \xordvalue~11 (
	.dataa(!dffe16),
	.datab(!dffe9),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~11 .extended_lut = "off";
defparam \xordvalue~11 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~11 .shared_arith = "off";

arriav_lcell_comb \xordvalue~12 (
	.dataa(!dffe16),
	.datab(!dffe10),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~12 .extended_lut = "off";
defparam \xordvalue~12 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~12 .shared_arith = "off";

endmodule

module nco_test_lpm_add_sub_4 (
	a_17,
	xordvalue_12,
	a_16,
	a_15,
	a_14,
	a_13,
	a_12,
	a_11,
	xordvalue_11,
	a_10,
	xordvalue_10,
	a_9,
	xordvalue_9,
	a_8,
	xordvalue_8,
	a_7,
	xordvalue_7,
	a_6,
	xordvalue_6,
	a_0,
	xordvalue_0,
	a_5,
	xordvalue_5,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	a_4,
	xordvalue_4,
	pipeline_dffe_17,
	pipeline_dffe_16,
	pipeline_dffe_15,
	pipeline_dffe_14,
	pipeline_dffe_13,
	pipeline_dffe_12,
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_12;
input 	a_16;
input 	a_15;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	xordvalue_11;
input 	a_10;
input 	xordvalue_10;
input 	a_9;
input 	xordvalue_9;
input 	a_8;
input 	xordvalue_8;
input 	a_7;
input 	xordvalue_7;
input 	a_6;
input 	xordvalue_6;
input 	a_0;
input 	xordvalue_0;
input 	a_5;
input 	xordvalue_5;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
input 	a_4;
input 	xordvalue_4;
output 	pipeline_dffe_17;
output 	pipeline_dffe_16;
output 	pipeline_dffe_15;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_add_sub_0qg_2 auto_generated(
	.a_17(a_17),
	.xordvalue_12(xordvalue_12),
	.a_16(a_16),
	.a_15(a_15),
	.a_14(a_14),
	.a_13(a_13),
	.a_12(a_12),
	.a_11(a_11),
	.xordvalue_11(xordvalue_11),
	.a_10(a_10),
	.xordvalue_10(xordvalue_10),
	.a_9(a_9),
	.xordvalue_9(xordvalue_9),
	.a_8(a_8),
	.xordvalue_8(xordvalue_8),
	.a_7(a_7),
	.xordvalue_7(xordvalue_7),
	.a_6(a_6),
	.xordvalue_6(xordvalue_6),
	.a_0(a_0),
	.xordvalue_0(xordvalue_0),
	.a_5(a_5),
	.xordvalue_5(xordvalue_5),
	.a_1(a_1),
	.xordvalue_1(xordvalue_1),
	.a_2(a_2),
	.xordvalue_2(xordvalue_2),
	.a_3(a_3),
	.xordvalue_3(xordvalue_3),
	.a_4(a_4),
	.xordvalue_4(xordvalue_4),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module nco_test_add_sub_0qg_2 (
	a_17,
	xordvalue_12,
	a_16,
	a_15,
	a_14,
	a_13,
	a_12,
	a_11,
	xordvalue_11,
	a_10,
	xordvalue_10,
	a_9,
	xordvalue_9,
	a_8,
	xordvalue_8,
	a_7,
	xordvalue_7,
	a_6,
	xordvalue_6,
	a_0,
	xordvalue_0,
	a_5,
	xordvalue_5,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	a_4,
	xordvalue_4,
	pipeline_dffe_17,
	pipeline_dffe_16,
	pipeline_dffe_15,
	pipeline_dffe_14,
	pipeline_dffe_13,
	pipeline_dffe_12,
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_12;
input 	a_16;
input 	a_15;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	xordvalue_11;
input 	a_10;
input 	xordvalue_10;
input 	a_9;
input 	xordvalue_9;
input 	a_8;
input 	xordvalue_8;
input 	a_7;
input 	xordvalue_7;
input 	a_6;
input 	xordvalue_6;
input 	a_0;
input 	xordvalue_0;
input 	a_5;
input 	xordvalue_5;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
input 	a_4;
input 	xordvalue_4;
output 	pipeline_dffe_17;
output 	pipeline_dffe_16;
output 	pipeline_dffe_15;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \op_1~50 ;
wire \op_1~58 ;
wire \op_1~62 ;
wire \op_1~66 ;
wire \op_1~70 ;
wire \op_1~54 ;
wire \op_1~46 ;
wire \op_1~42 ;
wire \op_1~38 ;
wire \op_1~34 ;
wire \op_1~30 ;
wire \op_1~26 ;
wire \op_1~22 ;
wire \op_1~18 ;
wire \op_1~14 ;
wire \op_1~10 ;
wire \op_1~6 ;
wire \op_1~1_sumout ;
wire \op_1~5_sumout ;
wire \op_1~9_sumout ;
wire \op_1~13_sumout ;
wire \op_1~17_sumout ;
wire \op_1~21_sumout ;
wire \op_1~25_sumout ;
wire \op_1~29_sumout ;
wire \op_1~33_sumout ;
wire \op_1~37_sumout ;
wire \op_1~45_sumout ;
wire \op_1~41_sumout ;
wire \op_1~49_sumout ;
wire \op_1~57_sumout ;
wire \op_1~61_sumout ;
wire \op_1~65_sumout ;
wire \op_1~69_sumout ;
wire \op_1~53_sumout ;


dffeas \pipeline_dffe[17] (
	.clk(clock),
	.d(\op_1~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_17),
	.prn(vcc));
defparam \pipeline_dffe[17] .is_wysiwyg = "true";
defparam \pipeline_dffe[17] .power_up = "low";

dffeas \pipeline_dffe[16] (
	.clk(clock),
	.d(\op_1~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_16),
	.prn(vcc));
defparam \pipeline_dffe[16] .is_wysiwyg = "true";
defparam \pipeline_dffe[16] .power_up = "low";

dffeas \pipeline_dffe[15] (
	.clk(clock),
	.d(\op_1~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_15),
	.prn(vcc));
defparam \pipeline_dffe[15] .is_wysiwyg = "true";
defparam \pipeline_dffe[15] .power_up = "low";

dffeas \pipeline_dffe[14] (
	.clk(clock),
	.d(\op_1~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_14),
	.prn(vcc));
defparam \pipeline_dffe[14] .is_wysiwyg = "true";
defparam \pipeline_dffe[14] .power_up = "low";

dffeas \pipeline_dffe[13] (
	.clk(clock),
	.d(\op_1~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_13),
	.prn(vcc));
defparam \pipeline_dffe[13] .is_wysiwyg = "true";
defparam \pipeline_dffe[13] .power_up = "low";

dffeas \pipeline_dffe[12] (
	.clk(clock),
	.d(\op_1~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_12),
	.prn(vcc));
defparam \pipeline_dffe[12] .is_wysiwyg = "true";
defparam \pipeline_dffe[12] .power_up = "low";

dffeas \pipeline_dffe[11] (
	.clk(clock),
	.d(\op_1~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \pipeline_dffe[11] .is_wysiwyg = "true";
defparam \pipeline_dffe[11] .power_up = "low";

dffeas \pipeline_dffe[10] (
	.clk(clock),
	.d(\op_1~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \pipeline_dffe[10] .is_wysiwyg = "true";
defparam \pipeline_dffe[10] .power_up = "low";

dffeas \pipeline_dffe[9] (
	.clk(clock),
	.d(\op_1~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \pipeline_dffe[9] .is_wysiwyg = "true";
defparam \pipeline_dffe[9] .power_up = "low";

dffeas \pipeline_dffe[8] (
	.clk(clock),
	.d(\op_1~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \pipeline_dffe[8] .is_wysiwyg = "true";
defparam \pipeline_dffe[8] .power_up = "low";

dffeas \pipeline_dffe[6] (
	.clk(clock),
	.d(\op_1~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \pipeline_dffe[6] .is_wysiwyg = "true";
defparam \pipeline_dffe[6] .power_up = "low";

dffeas \pipeline_dffe[7] (
	.clk(clock),
	.d(\op_1~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \pipeline_dffe[7] .is_wysiwyg = "true";
defparam \pipeline_dffe[7] .power_up = "low";

dffeas \pipeline_dffe[0] (
	.clk(clock),
	.d(\op_1~49_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_0),
	.prn(vcc));
defparam \pipeline_dffe[0] .is_wysiwyg = "true";
defparam \pipeline_dffe[0] .power_up = "low";

dffeas \pipeline_dffe[1] (
	.clk(clock),
	.d(\op_1~57_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_1),
	.prn(vcc));
defparam \pipeline_dffe[1] .is_wysiwyg = "true";
defparam \pipeline_dffe[1] .power_up = "low";

dffeas \pipeline_dffe[2] (
	.clk(clock),
	.d(\op_1~61_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \pipeline_dffe[2] .is_wysiwyg = "true";
defparam \pipeline_dffe[2] .power_up = "low";

dffeas \pipeline_dffe[3] (
	.clk(clock),
	.d(\op_1~65_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \pipeline_dffe[3] .is_wysiwyg = "true";
defparam \pipeline_dffe[3] .power_up = "low";

dffeas \pipeline_dffe[4] (
	.clk(clock),
	.d(\op_1~69_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \pipeline_dffe[4] .is_wysiwyg = "true";
defparam \pipeline_dffe[4] .power_up = "low";

dffeas \pipeline_dffe[5] (
	.clk(clock),
	.d(\op_1~53_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \pipeline_dffe[5] .is_wysiwyg = "true";
defparam \pipeline_dffe[5] .power_up = "low";

arriav_lcell_comb \op_1~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~49_sumout ),
	.cout(\op_1~50 ),
	.shareout());
defparam \op_1~49 .extended_lut = "off";
defparam \op_1~49 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~49 .shared_arith = "off";

arriav_lcell_comb \op_1~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_1),
	.datag(gnd),
	.cin(\op_1~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~57_sumout ),
	.cout(\op_1~58 ),
	.shareout());
defparam \op_1~57 .extended_lut = "off";
defparam \op_1~57 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~57 .shared_arith = "off";

arriav_lcell_comb \op_1~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_2),
	.datag(gnd),
	.cin(\op_1~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~61_sumout ),
	.cout(\op_1~62 ),
	.shareout());
defparam \op_1~61 .extended_lut = "off";
defparam \op_1~61 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~61 .shared_arith = "off";

arriav_lcell_comb \op_1~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_3),
	.datag(gnd),
	.cin(\op_1~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~65_sumout ),
	.cout(\op_1~66 ),
	.shareout());
defparam \op_1~65 .extended_lut = "off";
defparam \op_1~65 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~65 .shared_arith = "off";

arriav_lcell_comb \op_1~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_4),
	.datag(gnd),
	.cin(\op_1~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~69_sumout ),
	.cout(\op_1~70 ),
	.shareout());
defparam \op_1~69 .extended_lut = "off";
defparam \op_1~69 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~69 .shared_arith = "off";

arriav_lcell_comb \op_1~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_5),
	.datag(gnd),
	.cin(\op_1~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~53_sumout ),
	.cout(\op_1~54 ),
	.shareout());
defparam \op_1~53 .extended_lut = "off";
defparam \op_1~53 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~53 .shared_arith = "off";

arriav_lcell_comb \op_1~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_6),
	.datag(gnd),
	.cin(\op_1~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~45_sumout ),
	.cout(\op_1~46 ),
	.shareout());
defparam \op_1~45 .extended_lut = "off";
defparam \op_1~45 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~45 .shared_arith = "off";

arriav_lcell_comb \op_1~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_7),
	.datag(gnd),
	.cin(\op_1~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~41_sumout ),
	.cout(\op_1~42 ),
	.shareout());
defparam \op_1~41 .extended_lut = "off";
defparam \op_1~41 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~41 .shared_arith = "off";

arriav_lcell_comb \op_1~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_8),
	.datag(gnd),
	.cin(\op_1~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~37_sumout ),
	.cout(\op_1~38 ),
	.shareout());
defparam \op_1~37 .extended_lut = "off";
defparam \op_1~37 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~37 .shared_arith = "off";

arriav_lcell_comb \op_1~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_9),
	.datag(gnd),
	.cin(\op_1~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~33_sumout ),
	.cout(\op_1~34 ),
	.shareout());
defparam \op_1~33 .extended_lut = "off";
defparam \op_1~33 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~33 .shared_arith = "off";

arriav_lcell_comb \op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~29_sumout ),
	.cout(\op_1~30 ),
	.shareout());
defparam \op_1~29 .extended_lut = "off";
defparam \op_1~29 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~29 .shared_arith = "off";

arriav_lcell_comb \op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_11),
	.datag(gnd),
	.cin(\op_1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~25_sumout ),
	.cout(\op_1~26 ),
	.shareout());
defparam \op_1~25 .extended_lut = "off";
defparam \op_1~25 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~25 .shared_arith = "off";

arriav_lcell_comb \op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_12),
	.datag(gnd),
	.cin(\op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~21_sumout ),
	.cout(\op_1~22 ),
	.shareout());
defparam \op_1~21 .extended_lut = "off";
defparam \op_1~21 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~21 .shared_arith = "off";

arriav_lcell_comb \op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_12),
	.datag(gnd),
	.cin(\op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~17_sumout ),
	.cout(\op_1~18 ),
	.shareout());
defparam \op_1~17 .extended_lut = "off";
defparam \op_1~17 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~17 .shared_arith = "off";

arriav_lcell_comb \op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_12),
	.datag(gnd),
	.cin(\op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~13_sumout ),
	.cout(\op_1~14 ),
	.shareout());
defparam \op_1~13 .extended_lut = "off";
defparam \op_1~13 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~13 .shared_arith = "off";

arriav_lcell_comb \op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_12),
	.datag(gnd),
	.cin(\op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~9_sumout ),
	.cout(\op_1~10 ),
	.shareout());
defparam \op_1~9 .extended_lut = "off";
defparam \op_1~9 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~9 .shared_arith = "off";

arriav_lcell_comb \op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_16),
	.datae(gnd),
	.dataf(!xordvalue_12),
	.datag(gnd),
	.cin(\op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~5_sumout ),
	.cout(\op_1~6 ),
	.shareout());
defparam \op_1~5 .extended_lut = "off";
defparam \op_1~5 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~5 .shared_arith = "off";

arriav_lcell_comb \op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_17),
	.datae(gnd),
	.dataf(!xordvalue_12),
	.datag(gnd),
	.cin(\op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~1_sumout ),
	.cout(),
	.shareout());
defparam \op_1~1 .extended_lut = "off";
defparam \op_1~1 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~1 .shared_arith = "off";

endmodule

module nco_test_cordic_axor_1p_lpm_3 (
	sin_o_0,
	pipeline_dffe_17,
	pipeline_dffe_16,
	dffe16,
	pipeline_dffe_15,
	pipeline_dffe_171,
	dffe18,
	pipeline_dffe_14,
	pipeline_dffe_13,
	dffe17,
	pipeline_dffe_161,
	pipeline_dffe_12,
	dffe161,
	pipeline_dffe_151,
	pipeline_dffe_11,
	dffe15,
	pipeline_dffe_141,
	pipeline_dffe_10,
	dffe14,
	pipeline_dffe_131,
	pipeline_dffe_9,
	dffe13,
	pipeline_dffe_121,
	pipeline_dffe_8,
	dffe12,
	pipeline_dffe_7,
	pipeline_dffe_111,
	pipeline_dffe_0,
	dffe11,
	pipeline_dffe_101,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	dffe10,
	pipeline_dffe_91,
	dffe9,
	pipeline_dffe_81,
	dffe7,
	dffe8,
	pipeline_dffe_61,
	pipeline_dffe_71,
	pipeline_dffe_01,
	pipeline_dffe_18,
	pipeline_dffe_21,
	pipeline_dffe_31,
	pipeline_dffe_41,
	pipeline_dffe_51,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	sin_o_0;
output 	pipeline_dffe_17;
output 	pipeline_dffe_16;
input 	dffe16;
output 	pipeline_dffe_15;
input 	pipeline_dffe_171;
input 	dffe18;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
input 	dffe17;
input 	pipeline_dffe_161;
output 	pipeline_dffe_12;
input 	dffe161;
input 	pipeline_dffe_151;
output 	pipeline_dffe_11;
input 	dffe15;
input 	pipeline_dffe_141;
output 	pipeline_dffe_10;
input 	dffe14;
input 	pipeline_dffe_131;
output 	pipeline_dffe_9;
input 	dffe13;
input 	pipeline_dffe_121;
output 	pipeline_dffe_8;
input 	dffe12;
output 	pipeline_dffe_7;
input 	pipeline_dffe_111;
output 	pipeline_dffe_0;
input 	dffe11;
input 	pipeline_dffe_101;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
input 	dffe10;
input 	pipeline_dffe_91;
input 	dffe9;
input 	pipeline_dffe_81;
input 	dffe7;
input 	dffe8;
input 	pipeline_dffe_61;
input 	pipeline_dffe_71;
input 	pipeline_dffe_01;
input 	pipeline_dffe_18;
input 	pipeline_dffe_21;
input 	pipeline_dffe_31;
input 	pipeline_dffe_41;
input 	pipeline_dffe_51;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[17]~q ;
wire \xordvalue[11]~q ;
wire \Add0~1_sumout ;
wire \a[16]~q ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \a[15]~q ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \a[14]~q ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \a[13]~q ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \a[12]~q ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \a[11]~q ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \a[10]~q ;
wire \xordvalue[10]~q ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \a[9]~q ;
wire \xordvalue[9]~q ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \a[8]~q ;
wire \xordvalue[8]~q ;
wire \a[7]~q ;
wire \xordvalue[7]~q ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \a[0]~q ;
wire \xordvalue[0]~q ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \a[6]~q ;
wire \xordvalue[6]~q ;
wire \a[1]~q ;
wire \xordvalue[1]~q ;
wire \a[2]~q ;
wire \xordvalue[2]~q ;
wire \a[3]~q ;
wire \xordvalue[3]~q ;
wire \a[4]~q ;
wire \xordvalue[4]~q ;
wire \a[5]~q ;
wire \xordvalue[5]~q ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~65_sumout ;
wire \Add0~66 ;
wire \Add0~69_sumout ;
wire \Add0~70 ;
wire \xordvalue~0_combout ;
wire \xordvalue~1_combout ;
wire \xordvalue~2_combout ;
wire \xordvalue~3_combout ;
wire \xordvalue~4_combout ;
wire \xordvalue~5_combout ;
wire \xordvalue~6_combout ;
wire \xordvalue~7_combout ;
wire \xordvalue~8_combout ;
wire \xordvalue~9_combout ;
wire \xordvalue~10_combout ;
wire \xordvalue~11_combout ;


nco_test_lpm_add_sub_5 u0(
	.a_17(\a[17]~q ),
	.xordvalue_11(\xordvalue[11]~q ),
	.a_16(\a[16]~q ),
	.a_15(\a[15]~q ),
	.a_14(\a[14]~q ),
	.a_13(\a[13]~q ),
	.a_12(\a[12]~q ),
	.a_11(\a[11]~q ),
	.a_10(\a[10]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.a_9(\a[9]~q ),
	.xordvalue_9(\xordvalue[9]~q ),
	.a_8(\a[8]~q ),
	.xordvalue_8(\xordvalue[8]~q ),
	.a_7(\a[7]~q ),
	.xordvalue_7(\xordvalue[7]~q ),
	.a_0(\a[0]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_6(\a[6]~q ),
	.xordvalue_6(\xordvalue[6]~q ),
	.a_1(\a[1]~q ),
	.xordvalue_1(\xordvalue[1]~q ),
	.a_2(\a[2]~q ),
	.xordvalue_2(\xordvalue[2]~q ),
	.a_3(\a[3]~q ),
	.xordvalue_3(\xordvalue[3]~q ),
	.a_4(\a[4]~q ),
	.xordvalue_4(\xordvalue[4]~q ),
	.a_5(\a[5]~q ),
	.xordvalue_5(\xordvalue[5]~q ),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[17] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[17]~q ),
	.prn(vcc));
defparam \a[17] .is_wysiwyg = "true";
defparam \a[17] .power_up = "low";

dffeas \xordvalue[11] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[11]~q ),
	.prn(vcc));
defparam \xordvalue[11] .is_wysiwyg = "true";
defparam \xordvalue[11] .power_up = "low";

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_171),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h00000000000000FF;
defparam \Add0~1 .shared_arith = "off";

dffeas \a[16] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[16]~q ),
	.prn(vcc));
defparam \a[16] .is_wysiwyg = "true";
defparam \a[16] .power_up = "low";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h00000000000000FF;
defparam \Add0~5 .shared_arith = "off";

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h00000000000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h00000000000000FF;
defparam \Add0~13 .shared_arith = "off";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h00000000000000FF;
defparam \Add0~17 .shared_arith = "off";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h00000000000000FF;
defparam \Add0~21 .shared_arith = "off";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h00000000000000FF;
defparam \Add0~25 .shared_arith = "off";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(\xordvalue~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h00000000000000FF;
defparam \Add0~29 .shared_arith = "off";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \xordvalue[9] (
	.clk(clk),
	.d(\xordvalue~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[9]~q ),
	.prn(vcc));
defparam \xordvalue[9] .is_wysiwyg = "true";
defparam \xordvalue[9] .power_up = "low";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h00000000000000FF;
defparam \Add0~33 .shared_arith = "off";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \xordvalue[8] (
	.clk(clk),
	.d(\xordvalue~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[8]~q ),
	.prn(vcc));
defparam \xordvalue[8] .is_wysiwyg = "true";
defparam \xordvalue[8] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \xordvalue[7] (
	.clk(clk),
	.d(\xordvalue~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[7]~q ),
	.prn(vcc));
defparam \xordvalue[7] .is_wysiwyg = "true";
defparam \xordvalue[7] .power_up = "low";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h00000000000000FF;
defparam \Add0~37 .shared_arith = "off";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h00000000000000FF;
defparam \Add0~41 .shared_arith = "off";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \xordvalue[6] (
	.clk(clk),
	.d(\xordvalue~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[6]~q ),
	.prn(vcc));
defparam \xordvalue[6] .is_wysiwyg = "true";
defparam \xordvalue[6] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \xordvalue[1] (
	.clk(clk),
	.d(\xordvalue~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[1]~q ),
	.prn(vcc));
defparam \xordvalue[1] .is_wysiwyg = "true";
defparam \xordvalue[1] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \xordvalue[2] (
	.clk(clk),
	.d(\xordvalue~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[2]~q ),
	.prn(vcc));
defparam \xordvalue[2] .is_wysiwyg = "true";
defparam \xordvalue[2] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \xordvalue[3] (
	.clk(clk),
	.d(\xordvalue~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[3]~q ),
	.prn(vcc));
defparam \xordvalue[3] .is_wysiwyg = "true";
defparam \xordvalue[3] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \xordvalue[4] (
	.clk(clk),
	.d(\xordvalue~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[4]~q ),
	.prn(vcc));
defparam \xordvalue[4] .is_wysiwyg = "true";
defparam \xordvalue[4] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \xordvalue[5] (
	.clk(clk),
	.d(\xordvalue~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[5]~q ),
	.prn(vcc));
defparam \xordvalue[5] .is_wysiwyg = "true";
defparam \xordvalue[5] .power_up = "low";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe16),
	.datae(gnd),
	.dataf(!pipeline_dffe_01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~45 .shared_arith = "off";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout());
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h00000000000000FF;
defparam \Add0~49 .shared_arith = "off";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_18),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout());
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h00000000000000FF;
defparam \Add0~53 .shared_arith = "off";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout());
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h00000000000000FF;
defparam \Add0~57 .shared_arith = "off";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout());
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h00000000000000FF;
defparam \Add0~61 .shared_arith = "off";

arriav_lcell_comb \Add0~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~65_sumout ),
	.cout(\Add0~66 ),
	.shareout());
defparam \Add0~65 .extended_lut = "off";
defparam \Add0~65 .lut_mask = 64'h00000000000000FF;
defparam \Add0~65 .shared_arith = "off";

arriav_lcell_comb \Add0~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~69_sumout ),
	.cout(\Add0~70 ),
	.shareout());
defparam \Add0~69 .extended_lut = "off";
defparam \Add0~69 .lut_mask = 64'h00000000000000FF;
defparam \Add0~69 .shared_arith = "off";

arriav_lcell_comb \xordvalue~0 (
	.dataa(!dffe18),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

arriav_lcell_comb \xordvalue~1 (
	.dataa(!dffe17),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~1 .extended_lut = "off";
defparam \xordvalue~1 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~1 .shared_arith = "off";

arriav_lcell_comb \xordvalue~2 (
	.dataa(!dffe161),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~2 .extended_lut = "off";
defparam \xordvalue~2 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~2 .shared_arith = "off";

arriav_lcell_comb \xordvalue~3 (
	.dataa(!dffe15),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~3 .extended_lut = "off";
defparam \xordvalue~3 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~3 .shared_arith = "off";

arriav_lcell_comb \xordvalue~4 (
	.dataa(!dffe14),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~4 .extended_lut = "off";
defparam \xordvalue~4 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~4 .shared_arith = "off";

arriav_lcell_comb \xordvalue~5 (
	.dataa(!dffe7),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~5 .extended_lut = "off";
defparam \xordvalue~5 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~5 .shared_arith = "off";

arriav_lcell_comb \xordvalue~6 (
	.dataa(!dffe13),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~6 .extended_lut = "off";
defparam \xordvalue~6 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~6 .shared_arith = "off";

arriav_lcell_comb \xordvalue~7 (
	.dataa(!dffe8),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~7 .extended_lut = "off";
defparam \xordvalue~7 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~7 .shared_arith = "off";

arriav_lcell_comb \xordvalue~8 (
	.dataa(!dffe9),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~8 .extended_lut = "off";
defparam \xordvalue~8 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~8 .shared_arith = "off";

arriav_lcell_comb \xordvalue~9 (
	.dataa(!dffe10),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~9 .extended_lut = "off";
defparam \xordvalue~9 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~9 .shared_arith = "off";

arriav_lcell_comb \xordvalue~10 (
	.dataa(!dffe11),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~10 .extended_lut = "off";
defparam \xordvalue~10 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~10 .shared_arith = "off";

arriav_lcell_comb \xordvalue~11 (
	.dataa(!dffe12),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~11 .extended_lut = "off";
defparam \xordvalue~11 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~11 .shared_arith = "off";

endmodule

module nco_test_lpm_add_sub_5 (
	a_17,
	xordvalue_11,
	a_16,
	a_15,
	a_14,
	a_13,
	a_12,
	a_11,
	a_10,
	xordvalue_10,
	a_9,
	xordvalue_9,
	a_8,
	xordvalue_8,
	a_7,
	xordvalue_7,
	a_0,
	xordvalue_0,
	a_6,
	xordvalue_6,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	a_4,
	xordvalue_4,
	a_5,
	xordvalue_5,
	pipeline_dffe_17,
	pipeline_dffe_16,
	pipeline_dffe_15,
	pipeline_dffe_14,
	pipeline_dffe_13,
	pipeline_dffe_12,
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_7,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_11;
input 	a_16;
input 	a_15;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_10;
input 	xordvalue_10;
input 	a_9;
input 	xordvalue_9;
input 	a_8;
input 	xordvalue_8;
input 	a_7;
input 	xordvalue_7;
input 	a_0;
input 	xordvalue_0;
input 	a_6;
input 	xordvalue_6;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
input 	a_4;
input 	xordvalue_4;
input 	a_5;
input 	xordvalue_5;
output 	pipeline_dffe_17;
output 	pipeline_dffe_16;
output 	pipeline_dffe_15;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_7;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_add_sub_0qg_3 auto_generated(
	.a_17(a_17),
	.xordvalue_11(xordvalue_11),
	.a_16(a_16),
	.a_15(a_15),
	.a_14(a_14),
	.a_13(a_13),
	.a_12(a_12),
	.a_11(a_11),
	.a_10(a_10),
	.xordvalue_10(xordvalue_10),
	.a_9(a_9),
	.xordvalue_9(xordvalue_9),
	.a_8(a_8),
	.xordvalue_8(xordvalue_8),
	.a_7(a_7),
	.xordvalue_7(xordvalue_7),
	.a_0(a_0),
	.xordvalue_0(xordvalue_0),
	.a_6(a_6),
	.xordvalue_6(xordvalue_6),
	.a_1(a_1),
	.xordvalue_1(xordvalue_1),
	.a_2(a_2),
	.xordvalue_2(xordvalue_2),
	.a_3(a_3),
	.xordvalue_3(xordvalue_3),
	.a_4(a_4),
	.xordvalue_4(xordvalue_4),
	.a_5(a_5),
	.xordvalue_5(xordvalue_5),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module nco_test_add_sub_0qg_3 (
	a_17,
	xordvalue_11,
	a_16,
	a_15,
	a_14,
	a_13,
	a_12,
	a_11,
	a_10,
	xordvalue_10,
	a_9,
	xordvalue_9,
	a_8,
	xordvalue_8,
	a_7,
	xordvalue_7,
	a_0,
	xordvalue_0,
	a_6,
	xordvalue_6,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	a_4,
	xordvalue_4,
	a_5,
	xordvalue_5,
	pipeline_dffe_17,
	pipeline_dffe_16,
	pipeline_dffe_15,
	pipeline_dffe_14,
	pipeline_dffe_13,
	pipeline_dffe_12,
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_7,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_11;
input 	a_16;
input 	a_15;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_10;
input 	xordvalue_10;
input 	a_9;
input 	xordvalue_9;
input 	a_8;
input 	xordvalue_8;
input 	a_7;
input 	xordvalue_7;
input 	a_0;
input 	xordvalue_0;
input 	a_6;
input 	xordvalue_6;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
input 	a_4;
input 	xordvalue_4;
input 	a_5;
input 	xordvalue_5;
output 	pipeline_dffe_17;
output 	pipeline_dffe_16;
output 	pipeline_dffe_15;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_7;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \op_1~46 ;
wire \op_1~54 ;
wire \op_1~58 ;
wire \op_1~62 ;
wire \op_1~66 ;
wire \op_1~70 ;
wire \op_1~50 ;
wire \op_1~42 ;
wire \op_1~38 ;
wire \op_1~34 ;
wire \op_1~30 ;
wire \op_1~26 ;
wire \op_1~22 ;
wire \op_1~18 ;
wire \op_1~14 ;
wire \op_1~10 ;
wire \op_1~6 ;
wire \op_1~1_sumout ;
wire \op_1~5_sumout ;
wire \op_1~9_sumout ;
wire \op_1~13_sumout ;
wire \op_1~17_sumout ;
wire \op_1~21_sumout ;
wire \op_1~25_sumout ;
wire \op_1~29_sumout ;
wire \op_1~33_sumout ;
wire \op_1~37_sumout ;
wire \op_1~41_sumout ;
wire \op_1~45_sumout ;
wire \op_1~53_sumout ;
wire \op_1~57_sumout ;
wire \op_1~61_sumout ;
wire \op_1~65_sumout ;
wire \op_1~69_sumout ;
wire \op_1~49_sumout ;


dffeas \pipeline_dffe[17] (
	.clk(clock),
	.d(\op_1~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_17),
	.prn(vcc));
defparam \pipeline_dffe[17] .is_wysiwyg = "true";
defparam \pipeline_dffe[17] .power_up = "low";

dffeas \pipeline_dffe[16] (
	.clk(clock),
	.d(\op_1~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_16),
	.prn(vcc));
defparam \pipeline_dffe[16] .is_wysiwyg = "true";
defparam \pipeline_dffe[16] .power_up = "low";

dffeas \pipeline_dffe[15] (
	.clk(clock),
	.d(\op_1~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_15),
	.prn(vcc));
defparam \pipeline_dffe[15] .is_wysiwyg = "true";
defparam \pipeline_dffe[15] .power_up = "low";

dffeas \pipeline_dffe[14] (
	.clk(clock),
	.d(\op_1~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_14),
	.prn(vcc));
defparam \pipeline_dffe[14] .is_wysiwyg = "true";
defparam \pipeline_dffe[14] .power_up = "low";

dffeas \pipeline_dffe[13] (
	.clk(clock),
	.d(\op_1~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_13),
	.prn(vcc));
defparam \pipeline_dffe[13] .is_wysiwyg = "true";
defparam \pipeline_dffe[13] .power_up = "low";

dffeas \pipeline_dffe[12] (
	.clk(clock),
	.d(\op_1~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_12),
	.prn(vcc));
defparam \pipeline_dffe[12] .is_wysiwyg = "true";
defparam \pipeline_dffe[12] .power_up = "low";

dffeas \pipeline_dffe[11] (
	.clk(clock),
	.d(\op_1~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \pipeline_dffe[11] .is_wysiwyg = "true";
defparam \pipeline_dffe[11] .power_up = "low";

dffeas \pipeline_dffe[10] (
	.clk(clock),
	.d(\op_1~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \pipeline_dffe[10] .is_wysiwyg = "true";
defparam \pipeline_dffe[10] .power_up = "low";

dffeas \pipeline_dffe[9] (
	.clk(clock),
	.d(\op_1~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \pipeline_dffe[9] .is_wysiwyg = "true";
defparam \pipeline_dffe[9] .power_up = "low";

dffeas \pipeline_dffe[8] (
	.clk(clock),
	.d(\op_1~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \pipeline_dffe[8] .is_wysiwyg = "true";
defparam \pipeline_dffe[8] .power_up = "low";

dffeas \pipeline_dffe[7] (
	.clk(clock),
	.d(\op_1~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \pipeline_dffe[7] .is_wysiwyg = "true";
defparam \pipeline_dffe[7] .power_up = "low";

dffeas \pipeline_dffe[0] (
	.clk(clock),
	.d(\op_1~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_0),
	.prn(vcc));
defparam \pipeline_dffe[0] .is_wysiwyg = "true";
defparam \pipeline_dffe[0] .power_up = "low";

dffeas \pipeline_dffe[1] (
	.clk(clock),
	.d(\op_1~53_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_1),
	.prn(vcc));
defparam \pipeline_dffe[1] .is_wysiwyg = "true";
defparam \pipeline_dffe[1] .power_up = "low";

dffeas \pipeline_dffe[2] (
	.clk(clock),
	.d(\op_1~57_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \pipeline_dffe[2] .is_wysiwyg = "true";
defparam \pipeline_dffe[2] .power_up = "low";

dffeas \pipeline_dffe[3] (
	.clk(clock),
	.d(\op_1~61_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \pipeline_dffe[3] .is_wysiwyg = "true";
defparam \pipeline_dffe[3] .power_up = "low";

dffeas \pipeline_dffe[4] (
	.clk(clock),
	.d(\op_1~65_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \pipeline_dffe[4] .is_wysiwyg = "true";
defparam \pipeline_dffe[4] .power_up = "low";

dffeas \pipeline_dffe[5] (
	.clk(clock),
	.d(\op_1~69_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \pipeline_dffe[5] .is_wysiwyg = "true";
defparam \pipeline_dffe[5] .power_up = "low";

dffeas \pipeline_dffe[6] (
	.clk(clock),
	.d(\op_1~49_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \pipeline_dffe[6] .is_wysiwyg = "true";
defparam \pipeline_dffe[6] .power_up = "low";

arriav_lcell_comb \op_1~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~45_sumout ),
	.cout(\op_1~46 ),
	.shareout());
defparam \op_1~45 .extended_lut = "off";
defparam \op_1~45 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~45 .shared_arith = "off";

arriav_lcell_comb \op_1~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_1),
	.datag(gnd),
	.cin(\op_1~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~53_sumout ),
	.cout(\op_1~54 ),
	.shareout());
defparam \op_1~53 .extended_lut = "off";
defparam \op_1~53 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~53 .shared_arith = "off";

arriav_lcell_comb \op_1~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_2),
	.datag(gnd),
	.cin(\op_1~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~57_sumout ),
	.cout(\op_1~58 ),
	.shareout());
defparam \op_1~57 .extended_lut = "off";
defparam \op_1~57 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~57 .shared_arith = "off";

arriav_lcell_comb \op_1~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_3),
	.datag(gnd),
	.cin(\op_1~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~61_sumout ),
	.cout(\op_1~62 ),
	.shareout());
defparam \op_1~61 .extended_lut = "off";
defparam \op_1~61 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~61 .shared_arith = "off";

arriav_lcell_comb \op_1~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_4),
	.datag(gnd),
	.cin(\op_1~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~65_sumout ),
	.cout(\op_1~66 ),
	.shareout());
defparam \op_1~65 .extended_lut = "off";
defparam \op_1~65 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~65 .shared_arith = "off";

arriav_lcell_comb \op_1~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_5),
	.datag(gnd),
	.cin(\op_1~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~69_sumout ),
	.cout(\op_1~70 ),
	.shareout());
defparam \op_1~69 .extended_lut = "off";
defparam \op_1~69 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~69 .shared_arith = "off";

arriav_lcell_comb \op_1~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_6),
	.datag(gnd),
	.cin(\op_1~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~49_sumout ),
	.cout(\op_1~50 ),
	.shareout());
defparam \op_1~49 .extended_lut = "off";
defparam \op_1~49 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~49 .shared_arith = "off";

arriav_lcell_comb \op_1~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_7),
	.datag(gnd),
	.cin(\op_1~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~41_sumout ),
	.cout(\op_1~42 ),
	.shareout());
defparam \op_1~41 .extended_lut = "off";
defparam \op_1~41 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~41 .shared_arith = "off";

arriav_lcell_comb \op_1~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_8),
	.datag(gnd),
	.cin(\op_1~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~37_sumout ),
	.cout(\op_1~38 ),
	.shareout());
defparam \op_1~37 .extended_lut = "off";
defparam \op_1~37 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~37 .shared_arith = "off";

arriav_lcell_comb \op_1~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_9),
	.datag(gnd),
	.cin(\op_1~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~33_sumout ),
	.cout(\op_1~34 ),
	.shareout());
defparam \op_1~33 .extended_lut = "off";
defparam \op_1~33 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~33 .shared_arith = "off";

arriav_lcell_comb \op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~29_sumout ),
	.cout(\op_1~30 ),
	.shareout());
defparam \op_1~29 .extended_lut = "off";
defparam \op_1~29 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~29 .shared_arith = "off";

arriav_lcell_comb \op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_11),
	.datag(gnd),
	.cin(\op_1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~25_sumout ),
	.cout(\op_1~26 ),
	.shareout());
defparam \op_1~25 .extended_lut = "off";
defparam \op_1~25 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~25 .shared_arith = "off";

arriav_lcell_comb \op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_11),
	.datag(gnd),
	.cin(\op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~21_sumout ),
	.cout(\op_1~22 ),
	.shareout());
defparam \op_1~21 .extended_lut = "off";
defparam \op_1~21 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~21 .shared_arith = "off";

arriav_lcell_comb \op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_11),
	.datag(gnd),
	.cin(\op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~17_sumout ),
	.cout(\op_1~18 ),
	.shareout());
defparam \op_1~17 .extended_lut = "off";
defparam \op_1~17 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~17 .shared_arith = "off";

arriav_lcell_comb \op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_11),
	.datag(gnd),
	.cin(\op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~13_sumout ),
	.cout(\op_1~14 ),
	.shareout());
defparam \op_1~13 .extended_lut = "off";
defparam \op_1~13 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~13 .shared_arith = "off";

arriav_lcell_comb \op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_11),
	.datag(gnd),
	.cin(\op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~9_sumout ),
	.cout(\op_1~10 ),
	.shareout());
defparam \op_1~9 .extended_lut = "off";
defparam \op_1~9 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~9 .shared_arith = "off";

arriav_lcell_comb \op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_16),
	.datae(gnd),
	.dataf(!xordvalue_11),
	.datag(gnd),
	.cin(\op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~5_sumout ),
	.cout(\op_1~6 ),
	.shareout());
defparam \op_1~5 .extended_lut = "off";
defparam \op_1~5 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~5 .shared_arith = "off";

arriav_lcell_comb \op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_17),
	.datae(gnd),
	.dataf(!xordvalue_11),
	.datag(gnd),
	.cin(\op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~1_sumout ),
	.cout(),
	.shareout());
defparam \op_1~1 .extended_lut = "off";
defparam \op_1~1 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~1 .shared_arith = "off";

endmodule

module nco_test_cordic_axor_1p_lpm_4 (
	sin_o_0,
	pipeline_dffe_17,
	pipeline_dffe_16,
	dffe16,
	dffe18,
	pipeline_dffe_15,
	pipeline_dffe_171,
	pipeline_dffe_14,
	pipeline_dffe_161,
	pipeline_dffe_13,
	dffe17,
	pipeline_dffe_151,
	pipeline_dffe_12,
	dffe161,
	pipeline_dffe_141,
	pipeline_dffe_11,
	dffe15,
	pipeline_dffe_131,
	pipeline_dffe_10,
	dffe14,
	pipeline_dffe_121,
	pipeline_dffe_8,
	pipeline_dffe_9,
	dffe13,
	pipeline_dffe_0,
	pipeline_dffe_111,
	dffe12,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_101,
	dffe11,
	pipeline_dffe_91,
	dffe10,
	dffe8,
	dffe9,
	pipeline_dffe_81,
	pipeline_dffe_71,
	pipeline_dffe_01,
	pipeline_dffe_18,
	pipeline_dffe_21,
	pipeline_dffe_31,
	pipeline_dffe_41,
	pipeline_dffe_51,
	pipeline_dffe_61,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	sin_o_0;
output 	pipeline_dffe_17;
output 	pipeline_dffe_16;
input 	dffe16;
input 	dffe18;
output 	pipeline_dffe_15;
input 	pipeline_dffe_171;
output 	pipeline_dffe_14;
input 	pipeline_dffe_161;
output 	pipeline_dffe_13;
input 	dffe17;
input 	pipeline_dffe_151;
output 	pipeline_dffe_12;
input 	dffe161;
input 	pipeline_dffe_141;
output 	pipeline_dffe_11;
input 	dffe15;
input 	pipeline_dffe_131;
output 	pipeline_dffe_10;
input 	dffe14;
input 	pipeline_dffe_121;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	dffe13;
output 	pipeline_dffe_0;
input 	pipeline_dffe_111;
input 	dffe12;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
input 	pipeline_dffe_101;
input 	dffe11;
input 	pipeline_dffe_91;
input 	dffe10;
input 	dffe8;
input 	dffe9;
input 	pipeline_dffe_81;
input 	pipeline_dffe_71;
input 	pipeline_dffe_01;
input 	pipeline_dffe_18;
input 	pipeline_dffe_21;
input 	pipeline_dffe_31;
input 	pipeline_dffe_41;
input 	pipeline_dffe_51;
input 	pipeline_dffe_61;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[17]~q ;
wire \xordvalue[10]~q ;
wire \Add0~1_sumout ;
wire \a[16]~q ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \a[15]~q ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \a[14]~q ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \a[13]~q ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \a[12]~q ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \a[11]~q ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \a[10]~q ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \a[9]~q ;
wire \xordvalue[9]~q ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \a[8]~q ;
wire \xordvalue[8]~q ;
wire \a[0]~q ;
wire \xordvalue[0]~q ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \a[7]~q ;
wire \xordvalue[7]~q ;
wire \a[1]~q ;
wire \xordvalue[1]~q ;
wire \a[2]~q ;
wire \xordvalue[2]~q ;
wire \a[3]~q ;
wire \xordvalue[3]~q ;
wire \a[4]~q ;
wire \xordvalue[4]~q ;
wire \a[5]~q ;
wire \xordvalue[5]~q ;
wire \a[6]~q ;
wire \xordvalue[6]~q ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~65_sumout ;
wire \Add0~66 ;
wire \Add0~69_sumout ;
wire \Add0~70 ;
wire \xordvalue~0_combout ;
wire \xordvalue~1_combout ;
wire \xordvalue~2_combout ;
wire \xordvalue~3_combout ;
wire \xordvalue~4_combout ;
wire \xordvalue~5_combout ;
wire \xordvalue~6_combout ;
wire \xordvalue~7_combout ;
wire \xordvalue~8_combout ;
wire \xordvalue~9_combout ;
wire \xordvalue~10_combout ;


nco_test_lpm_add_sub_6 u0(
	.a_17(\a[17]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.a_16(\a[16]~q ),
	.a_15(\a[15]~q ),
	.a_14(\a[14]~q ),
	.a_13(\a[13]~q ),
	.a_12(\a[12]~q ),
	.a_11(\a[11]~q ),
	.a_10(\a[10]~q ),
	.a_9(\a[9]~q ),
	.xordvalue_9(\xordvalue[9]~q ),
	.a_8(\a[8]~q ),
	.xordvalue_8(\xordvalue[8]~q ),
	.a_0(\a[0]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_7(\a[7]~q ),
	.xordvalue_7(\xordvalue[7]~q ),
	.a_1(\a[1]~q ),
	.xordvalue_1(\xordvalue[1]~q ),
	.a_2(\a[2]~q ),
	.xordvalue_2(\xordvalue[2]~q ),
	.a_3(\a[3]~q ),
	.xordvalue_3(\xordvalue[3]~q ),
	.a_4(\a[4]~q ),
	.xordvalue_4(\xordvalue[4]~q ),
	.a_5(\a[5]~q ),
	.xordvalue_5(\xordvalue[5]~q ),
	.a_6(\a[6]~q ),
	.xordvalue_6(\xordvalue[6]~q ),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[17] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[17]~q ),
	.prn(vcc));
defparam \a[17] .is_wysiwyg = "true";
defparam \a[17] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_171),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h00000000000000FF;
defparam \Add0~1 .shared_arith = "off";

dffeas \a[16] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[16]~q ),
	.prn(vcc));
defparam \a[16] .is_wysiwyg = "true";
defparam \a[16] .power_up = "low";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h00000000000000FF;
defparam \Add0~5 .shared_arith = "off";

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h00000000000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h00000000000000FF;
defparam \Add0~13 .shared_arith = "off";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h00000000000000FF;
defparam \Add0~17 .shared_arith = "off";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h00000000000000FF;
defparam \Add0~21 .shared_arith = "off";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h00000000000000FF;
defparam \Add0~25 .shared_arith = "off";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h00000000000000FF;
defparam \Add0~29 .shared_arith = "off";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \xordvalue[9] (
	.clk(clk),
	.d(\xordvalue~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[9]~q ),
	.prn(vcc));
defparam \xordvalue[9] .is_wysiwyg = "true";
defparam \xordvalue[9] .power_up = "low";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h00000000000000FF;
defparam \Add0~33 .shared_arith = "off";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \xordvalue[8] (
	.clk(clk),
	.d(\xordvalue~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[8]~q ),
	.prn(vcc));
defparam \xordvalue[8] .is_wysiwyg = "true";
defparam \xordvalue[8] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h00000000000000FF;
defparam \Add0~37 .shared_arith = "off";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \xordvalue[7] (
	.clk(clk),
	.d(\xordvalue~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[7]~q ),
	.prn(vcc));
defparam \xordvalue[7] .is_wysiwyg = "true";
defparam \xordvalue[7] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \xordvalue[1] (
	.clk(clk),
	.d(\xordvalue~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[1]~q ),
	.prn(vcc));
defparam \xordvalue[1] .is_wysiwyg = "true";
defparam \xordvalue[1] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \xordvalue[2] (
	.clk(clk),
	.d(\xordvalue~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[2]~q ),
	.prn(vcc));
defparam \xordvalue[2] .is_wysiwyg = "true";
defparam \xordvalue[2] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \xordvalue[3] (
	.clk(clk),
	.d(\xordvalue~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[3]~q ),
	.prn(vcc));
defparam \xordvalue[3] .is_wysiwyg = "true";
defparam \xordvalue[3] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \xordvalue[4] (
	.clk(clk),
	.d(\xordvalue~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[4]~q ),
	.prn(vcc));
defparam \xordvalue[4] .is_wysiwyg = "true";
defparam \xordvalue[4] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \xordvalue[5] (
	.clk(clk),
	.d(\xordvalue~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[5]~q ),
	.prn(vcc));
defparam \xordvalue[5] .is_wysiwyg = "true";
defparam \xordvalue[5] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \xordvalue[6] (
	.clk(clk),
	.d(\xordvalue~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[6]~q ),
	.prn(vcc));
defparam \xordvalue[6] .is_wysiwyg = "true";
defparam \xordvalue[6] .power_up = "low";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe16),
	.datae(gnd),
	.dataf(!pipeline_dffe_01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~41 .shared_arith = "off";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h00000000000000FF;
defparam \Add0~45 .shared_arith = "off";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_18),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout());
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h00000000000000FF;
defparam \Add0~49 .shared_arith = "off";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout());
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h00000000000000FF;
defparam \Add0~53 .shared_arith = "off";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout());
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h00000000000000FF;
defparam \Add0~57 .shared_arith = "off";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout());
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h00000000000000FF;
defparam \Add0~61 .shared_arith = "off";

arriav_lcell_comb \Add0~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~65_sumout ),
	.cout(\Add0~66 ),
	.shareout());
defparam \Add0~65 .extended_lut = "off";
defparam \Add0~65 .lut_mask = 64'h00000000000000FF;
defparam \Add0~65 .shared_arith = "off";

arriav_lcell_comb \Add0~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~69_sumout ),
	.cout(\Add0~70 ),
	.shareout());
defparam \Add0~69 .extended_lut = "off";
defparam \Add0~69 .lut_mask = 64'h00000000000000FF;
defparam \Add0~69 .shared_arith = "off";

arriav_lcell_comb \xordvalue~0 (
	.dataa(!dffe16),
	.datab(!dffe18),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

arriav_lcell_comb \xordvalue~1 (
	.dataa(!dffe16),
	.datab(!dffe17),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~1 .extended_lut = "off";
defparam \xordvalue~1 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~1 .shared_arith = "off";

arriav_lcell_comb \xordvalue~2 (
	.dataa(!dffe16),
	.datab(!dffe161),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~2 .extended_lut = "off";
defparam \xordvalue~2 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~2 .shared_arith = "off";

arriav_lcell_comb \xordvalue~3 (
	.dataa(!dffe16),
	.datab(!dffe8),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~3 .extended_lut = "off";
defparam \xordvalue~3 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~3 .shared_arith = "off";

arriav_lcell_comb \xordvalue~4 (
	.dataa(!dffe16),
	.datab(!dffe15),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~4 .extended_lut = "off";
defparam \xordvalue~4 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~4 .shared_arith = "off";

arriav_lcell_comb \xordvalue~5 (
	.dataa(!dffe16),
	.datab(!dffe9),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~5 .extended_lut = "off";
defparam \xordvalue~5 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~5 .shared_arith = "off";

arriav_lcell_comb \xordvalue~6 (
	.dataa(!dffe16),
	.datab(!dffe10),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~6 .extended_lut = "off";
defparam \xordvalue~6 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~6 .shared_arith = "off";

arriav_lcell_comb \xordvalue~7 (
	.dataa(!dffe16),
	.datab(!dffe11),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~7 .extended_lut = "off";
defparam \xordvalue~7 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~7 .shared_arith = "off";

arriav_lcell_comb \xordvalue~8 (
	.dataa(!dffe16),
	.datab(!dffe12),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~8 .extended_lut = "off";
defparam \xordvalue~8 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~8 .shared_arith = "off";

arriav_lcell_comb \xordvalue~9 (
	.dataa(!dffe16),
	.datab(!dffe13),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~9 .extended_lut = "off";
defparam \xordvalue~9 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~9 .shared_arith = "off";

arriav_lcell_comb \xordvalue~10 (
	.dataa(!dffe16),
	.datab(!dffe14),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~10 .extended_lut = "off";
defparam \xordvalue~10 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~10 .shared_arith = "off";

endmodule

module nco_test_lpm_add_sub_6 (
	a_17,
	xordvalue_10,
	a_16,
	a_15,
	a_14,
	a_13,
	a_12,
	a_11,
	a_10,
	a_9,
	xordvalue_9,
	a_8,
	xordvalue_8,
	a_0,
	xordvalue_0,
	a_7,
	xordvalue_7,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	a_4,
	xordvalue_4,
	a_5,
	xordvalue_5,
	a_6,
	xordvalue_6,
	pipeline_dffe_17,
	pipeline_dffe_16,
	pipeline_dffe_15,
	pipeline_dffe_14,
	pipeline_dffe_13,
	pipeline_dffe_12,
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_10;
input 	a_16;
input 	a_15;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_10;
input 	a_9;
input 	xordvalue_9;
input 	a_8;
input 	xordvalue_8;
input 	a_0;
input 	xordvalue_0;
input 	a_7;
input 	xordvalue_7;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
input 	a_4;
input 	xordvalue_4;
input 	a_5;
input 	xordvalue_5;
input 	a_6;
input 	xordvalue_6;
output 	pipeline_dffe_17;
output 	pipeline_dffe_16;
output 	pipeline_dffe_15;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_add_sub_0qg_4 auto_generated(
	.a_17(a_17),
	.xordvalue_10(xordvalue_10),
	.a_16(a_16),
	.a_15(a_15),
	.a_14(a_14),
	.a_13(a_13),
	.a_12(a_12),
	.a_11(a_11),
	.a_10(a_10),
	.a_9(a_9),
	.xordvalue_9(xordvalue_9),
	.a_8(a_8),
	.xordvalue_8(xordvalue_8),
	.a_0(a_0),
	.xordvalue_0(xordvalue_0),
	.a_7(a_7),
	.xordvalue_7(xordvalue_7),
	.a_1(a_1),
	.xordvalue_1(xordvalue_1),
	.a_2(a_2),
	.xordvalue_2(xordvalue_2),
	.a_3(a_3),
	.xordvalue_3(xordvalue_3),
	.a_4(a_4),
	.xordvalue_4(xordvalue_4),
	.a_5(a_5),
	.xordvalue_5(xordvalue_5),
	.a_6(a_6),
	.xordvalue_6(xordvalue_6),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module nco_test_add_sub_0qg_4 (
	a_17,
	xordvalue_10,
	a_16,
	a_15,
	a_14,
	a_13,
	a_12,
	a_11,
	a_10,
	a_9,
	xordvalue_9,
	a_8,
	xordvalue_8,
	a_0,
	xordvalue_0,
	a_7,
	xordvalue_7,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	a_4,
	xordvalue_4,
	a_5,
	xordvalue_5,
	a_6,
	xordvalue_6,
	pipeline_dffe_17,
	pipeline_dffe_16,
	pipeline_dffe_15,
	pipeline_dffe_14,
	pipeline_dffe_13,
	pipeline_dffe_12,
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_10;
input 	a_16;
input 	a_15;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_10;
input 	a_9;
input 	xordvalue_9;
input 	a_8;
input 	xordvalue_8;
input 	a_0;
input 	xordvalue_0;
input 	a_7;
input 	xordvalue_7;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
input 	a_4;
input 	xordvalue_4;
input 	a_5;
input 	xordvalue_5;
input 	a_6;
input 	xordvalue_6;
output 	pipeline_dffe_17;
output 	pipeline_dffe_16;
output 	pipeline_dffe_15;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \op_1~42 ;
wire \op_1~50 ;
wire \op_1~54 ;
wire \op_1~58 ;
wire \op_1~62 ;
wire \op_1~66 ;
wire \op_1~70 ;
wire \op_1~46 ;
wire \op_1~38 ;
wire \op_1~34 ;
wire \op_1~30 ;
wire \op_1~26 ;
wire \op_1~22 ;
wire \op_1~18 ;
wire \op_1~14 ;
wire \op_1~10 ;
wire \op_1~6 ;
wire \op_1~1_sumout ;
wire \op_1~5_sumout ;
wire \op_1~9_sumout ;
wire \op_1~13_sumout ;
wire \op_1~17_sumout ;
wire \op_1~21_sumout ;
wire \op_1~25_sumout ;
wire \op_1~29_sumout ;
wire \op_1~37_sumout ;
wire \op_1~33_sumout ;
wire \op_1~41_sumout ;
wire \op_1~49_sumout ;
wire \op_1~53_sumout ;
wire \op_1~57_sumout ;
wire \op_1~61_sumout ;
wire \op_1~65_sumout ;
wire \op_1~69_sumout ;
wire \op_1~45_sumout ;


dffeas \pipeline_dffe[17] (
	.clk(clock),
	.d(\op_1~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_17),
	.prn(vcc));
defparam \pipeline_dffe[17] .is_wysiwyg = "true";
defparam \pipeline_dffe[17] .power_up = "low";

dffeas \pipeline_dffe[16] (
	.clk(clock),
	.d(\op_1~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_16),
	.prn(vcc));
defparam \pipeline_dffe[16] .is_wysiwyg = "true";
defparam \pipeline_dffe[16] .power_up = "low";

dffeas \pipeline_dffe[15] (
	.clk(clock),
	.d(\op_1~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_15),
	.prn(vcc));
defparam \pipeline_dffe[15] .is_wysiwyg = "true";
defparam \pipeline_dffe[15] .power_up = "low";

dffeas \pipeline_dffe[14] (
	.clk(clock),
	.d(\op_1~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_14),
	.prn(vcc));
defparam \pipeline_dffe[14] .is_wysiwyg = "true";
defparam \pipeline_dffe[14] .power_up = "low";

dffeas \pipeline_dffe[13] (
	.clk(clock),
	.d(\op_1~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_13),
	.prn(vcc));
defparam \pipeline_dffe[13] .is_wysiwyg = "true";
defparam \pipeline_dffe[13] .power_up = "low";

dffeas \pipeline_dffe[12] (
	.clk(clock),
	.d(\op_1~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_12),
	.prn(vcc));
defparam \pipeline_dffe[12] .is_wysiwyg = "true";
defparam \pipeline_dffe[12] .power_up = "low";

dffeas \pipeline_dffe[11] (
	.clk(clock),
	.d(\op_1~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \pipeline_dffe[11] .is_wysiwyg = "true";
defparam \pipeline_dffe[11] .power_up = "low";

dffeas \pipeline_dffe[10] (
	.clk(clock),
	.d(\op_1~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \pipeline_dffe[10] .is_wysiwyg = "true";
defparam \pipeline_dffe[10] .power_up = "low";

dffeas \pipeline_dffe[8] (
	.clk(clock),
	.d(\op_1~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \pipeline_dffe[8] .is_wysiwyg = "true";
defparam \pipeline_dffe[8] .power_up = "low";

dffeas \pipeline_dffe[9] (
	.clk(clock),
	.d(\op_1~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \pipeline_dffe[9] .is_wysiwyg = "true";
defparam \pipeline_dffe[9] .power_up = "low";

dffeas \pipeline_dffe[0] (
	.clk(clock),
	.d(\op_1~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_0),
	.prn(vcc));
defparam \pipeline_dffe[0] .is_wysiwyg = "true";
defparam \pipeline_dffe[0] .power_up = "low";

dffeas \pipeline_dffe[1] (
	.clk(clock),
	.d(\op_1~49_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_1),
	.prn(vcc));
defparam \pipeline_dffe[1] .is_wysiwyg = "true";
defparam \pipeline_dffe[1] .power_up = "low";

dffeas \pipeline_dffe[2] (
	.clk(clock),
	.d(\op_1~53_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \pipeline_dffe[2] .is_wysiwyg = "true";
defparam \pipeline_dffe[2] .power_up = "low";

dffeas \pipeline_dffe[3] (
	.clk(clock),
	.d(\op_1~57_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \pipeline_dffe[3] .is_wysiwyg = "true";
defparam \pipeline_dffe[3] .power_up = "low";

dffeas \pipeline_dffe[4] (
	.clk(clock),
	.d(\op_1~61_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \pipeline_dffe[4] .is_wysiwyg = "true";
defparam \pipeline_dffe[4] .power_up = "low";

dffeas \pipeline_dffe[5] (
	.clk(clock),
	.d(\op_1~65_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \pipeline_dffe[5] .is_wysiwyg = "true";
defparam \pipeline_dffe[5] .power_up = "low";

dffeas \pipeline_dffe[6] (
	.clk(clock),
	.d(\op_1~69_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \pipeline_dffe[6] .is_wysiwyg = "true";
defparam \pipeline_dffe[6] .power_up = "low";

dffeas \pipeline_dffe[7] (
	.clk(clock),
	.d(\op_1~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \pipeline_dffe[7] .is_wysiwyg = "true";
defparam \pipeline_dffe[7] .power_up = "low";

arriav_lcell_comb \op_1~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~41_sumout ),
	.cout(\op_1~42 ),
	.shareout());
defparam \op_1~41 .extended_lut = "off";
defparam \op_1~41 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~41 .shared_arith = "off";

arriav_lcell_comb \op_1~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_1),
	.datag(gnd),
	.cin(\op_1~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~49_sumout ),
	.cout(\op_1~50 ),
	.shareout());
defparam \op_1~49 .extended_lut = "off";
defparam \op_1~49 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~49 .shared_arith = "off";

arriav_lcell_comb \op_1~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_2),
	.datag(gnd),
	.cin(\op_1~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~53_sumout ),
	.cout(\op_1~54 ),
	.shareout());
defparam \op_1~53 .extended_lut = "off";
defparam \op_1~53 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~53 .shared_arith = "off";

arriav_lcell_comb \op_1~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_3),
	.datag(gnd),
	.cin(\op_1~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~57_sumout ),
	.cout(\op_1~58 ),
	.shareout());
defparam \op_1~57 .extended_lut = "off";
defparam \op_1~57 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~57 .shared_arith = "off";

arriav_lcell_comb \op_1~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_4),
	.datag(gnd),
	.cin(\op_1~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~61_sumout ),
	.cout(\op_1~62 ),
	.shareout());
defparam \op_1~61 .extended_lut = "off";
defparam \op_1~61 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~61 .shared_arith = "off";

arriav_lcell_comb \op_1~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_5),
	.datag(gnd),
	.cin(\op_1~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~65_sumout ),
	.cout(\op_1~66 ),
	.shareout());
defparam \op_1~65 .extended_lut = "off";
defparam \op_1~65 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~65 .shared_arith = "off";

arriav_lcell_comb \op_1~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_6),
	.datag(gnd),
	.cin(\op_1~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~69_sumout ),
	.cout(\op_1~70 ),
	.shareout());
defparam \op_1~69 .extended_lut = "off";
defparam \op_1~69 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~69 .shared_arith = "off";

arriav_lcell_comb \op_1~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_7),
	.datag(gnd),
	.cin(\op_1~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~45_sumout ),
	.cout(\op_1~46 ),
	.shareout());
defparam \op_1~45 .extended_lut = "off";
defparam \op_1~45 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~45 .shared_arith = "off";

arriav_lcell_comb \op_1~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_8),
	.datag(gnd),
	.cin(\op_1~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~37_sumout ),
	.cout(\op_1~38 ),
	.shareout());
defparam \op_1~37 .extended_lut = "off";
defparam \op_1~37 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~37 .shared_arith = "off";

arriav_lcell_comb \op_1~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_9),
	.datag(gnd),
	.cin(\op_1~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~33_sumout ),
	.cout(\op_1~34 ),
	.shareout());
defparam \op_1~33 .extended_lut = "off";
defparam \op_1~33 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~33 .shared_arith = "off";

arriav_lcell_comb \op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~29_sumout ),
	.cout(\op_1~30 ),
	.shareout());
defparam \op_1~29 .extended_lut = "off";
defparam \op_1~29 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~29 .shared_arith = "off";

arriav_lcell_comb \op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~25_sumout ),
	.cout(\op_1~26 ),
	.shareout());
defparam \op_1~25 .extended_lut = "off";
defparam \op_1~25 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~25 .shared_arith = "off";

arriav_lcell_comb \op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~21_sumout ),
	.cout(\op_1~22 ),
	.shareout());
defparam \op_1~21 .extended_lut = "off";
defparam \op_1~21 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~21 .shared_arith = "off";

arriav_lcell_comb \op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~17_sumout ),
	.cout(\op_1~18 ),
	.shareout());
defparam \op_1~17 .extended_lut = "off";
defparam \op_1~17 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~17 .shared_arith = "off";

arriav_lcell_comb \op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~13_sumout ),
	.cout(\op_1~14 ),
	.shareout());
defparam \op_1~13 .extended_lut = "off";
defparam \op_1~13 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~13 .shared_arith = "off";

arriav_lcell_comb \op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~9_sumout ),
	.cout(\op_1~10 ),
	.shareout());
defparam \op_1~9 .extended_lut = "off";
defparam \op_1~9 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~9 .shared_arith = "off";

arriav_lcell_comb \op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_16),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~5_sumout ),
	.cout(\op_1~6 ),
	.shareout());
defparam \op_1~5 .extended_lut = "off";
defparam \op_1~5 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~5 .shared_arith = "off";

arriav_lcell_comb \op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_17),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~1_sumout ),
	.cout(),
	.shareout());
defparam \op_1~1 .extended_lut = "off";
defparam \op_1~1 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~1 .shared_arith = "off";

endmodule

module nco_test_cordic_axor_1p_lpm_5 (
	sin_o_0,
	pipeline_dffe_17,
	pipeline_dffe_16,
	dffe16,
	pipeline_dffe_15,
	pipeline_dffe_171,
	dffe18,
	pipeline_dffe_14,
	pipeline_dffe_13,
	dffe17,
	pipeline_dffe_161,
	pipeline_dffe_12,
	dffe161,
	pipeline_dffe_151,
	pipeline_dffe_11,
	dffe15,
	pipeline_dffe_141,
	pipeline_dffe_10,
	dffe14,
	pipeline_dffe_9,
	pipeline_dffe_131,
	pipeline_dffe_0,
	dffe13,
	pipeline_dffe_121,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	dffe12,
	pipeline_dffe_111,
	dffe11,
	pipeline_dffe_101,
	dffe9,
	dffe10,
	pipeline_dffe_81,
	pipeline_dffe_91,
	pipeline_dffe_01,
	pipeline_dffe_18,
	pipeline_dffe_21,
	pipeline_dffe_31,
	pipeline_dffe_41,
	pipeline_dffe_51,
	pipeline_dffe_61,
	pipeline_dffe_71,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	sin_o_0;
output 	pipeline_dffe_17;
output 	pipeline_dffe_16;
input 	dffe16;
output 	pipeline_dffe_15;
input 	pipeline_dffe_171;
input 	dffe18;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
input 	dffe17;
input 	pipeline_dffe_161;
output 	pipeline_dffe_12;
input 	dffe161;
input 	pipeline_dffe_151;
output 	pipeline_dffe_11;
input 	dffe15;
input 	pipeline_dffe_141;
output 	pipeline_dffe_10;
input 	dffe14;
output 	pipeline_dffe_9;
input 	pipeline_dffe_131;
output 	pipeline_dffe_0;
input 	dffe13;
input 	pipeline_dffe_121;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
input 	dffe12;
input 	pipeline_dffe_111;
input 	dffe11;
input 	pipeline_dffe_101;
input 	dffe9;
input 	dffe10;
input 	pipeline_dffe_81;
input 	pipeline_dffe_91;
input 	pipeline_dffe_01;
input 	pipeline_dffe_18;
input 	pipeline_dffe_21;
input 	pipeline_dffe_31;
input 	pipeline_dffe_41;
input 	pipeline_dffe_51;
input 	pipeline_dffe_61;
input 	pipeline_dffe_71;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[17]~q ;
wire \xordvalue[10]~q ;
wire \Add0~1_sumout ;
wire \a[16]~q ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \a[15]~q ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \a[14]~q ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \a[13]~q ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \a[12]~q ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \a[11]~q ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \a[10]~q ;
wire \a[9]~q ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \a[0]~q ;
wire \xordvalue[0]~q ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \a[8]~q ;
wire \xordvalue[8]~q ;
wire \a[1]~q ;
wire \xordvalue[1]~q ;
wire \a[2]~q ;
wire \xordvalue[2]~q ;
wire \a[3]~q ;
wire \xordvalue[3]~q ;
wire \a[4]~q ;
wire \xordvalue[4]~q ;
wire \a[5]~q ;
wire \xordvalue[5]~q ;
wire \a[6]~q ;
wire \xordvalue[6]~q ;
wire \a[7]~q ;
wire \xordvalue[7]~q ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~65_sumout ;
wire \Add0~66 ;
wire \Add0~69_sumout ;
wire \Add0~70 ;
wire \xordvalue~0_combout ;
wire \xordvalue~1_combout ;
wire \xordvalue~2_combout ;
wire \xordvalue~3_combout ;
wire \xordvalue~4_combout ;
wire \xordvalue~5_combout ;
wire \xordvalue~6_combout ;
wire \xordvalue~7_combout ;
wire \xordvalue~8_combout ;
wire \xordvalue~9_combout ;


nco_test_lpm_add_sub_7 u0(
	.a_17(\a[17]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.a_16(\a[16]~q ),
	.a_15(\a[15]~q ),
	.a_14(\a[14]~q ),
	.a_13(\a[13]~q ),
	.a_12(\a[12]~q ),
	.a_11(\a[11]~q ),
	.a_10(\a[10]~q ),
	.a_9(\a[9]~q ),
	.a_0(\a[0]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_8(\a[8]~q ),
	.xordvalue_8(\xordvalue[8]~q ),
	.a_1(\a[1]~q ),
	.xordvalue_1(\xordvalue[1]~q ),
	.a_2(\a[2]~q ),
	.xordvalue_2(\xordvalue[2]~q ),
	.a_3(\a[3]~q ),
	.xordvalue_3(\xordvalue[3]~q ),
	.a_4(\a[4]~q ),
	.xordvalue_4(\xordvalue[4]~q ),
	.a_5(\a[5]~q ),
	.xordvalue_5(\xordvalue[5]~q ),
	.a_6(\a[6]~q ),
	.xordvalue_6(\xordvalue[6]~q ),
	.a_7(\a[7]~q ),
	.xordvalue_7(\xordvalue[7]~q ),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[17] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[17]~q ),
	.prn(vcc));
defparam \a[17] .is_wysiwyg = "true";
defparam \a[17] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_171),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h00000000000000FF;
defparam \Add0~1 .shared_arith = "off";

dffeas \a[16] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[16]~q ),
	.prn(vcc));
defparam \a[16] .is_wysiwyg = "true";
defparam \a[16] .power_up = "low";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h00000000000000FF;
defparam \Add0~5 .shared_arith = "off";

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h00000000000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h00000000000000FF;
defparam \Add0~13 .shared_arith = "off";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h00000000000000FF;
defparam \Add0~17 .shared_arith = "off";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h00000000000000FF;
defparam \Add0~21 .shared_arith = "off";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h00000000000000FF;
defparam \Add0~25 .shared_arith = "off";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h00000000000000FF;
defparam \Add0~29 .shared_arith = "off";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h00000000000000FF;
defparam \Add0~33 .shared_arith = "off";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \xordvalue[8] (
	.clk(clk),
	.d(\xordvalue~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[8]~q ),
	.prn(vcc));
defparam \xordvalue[8] .is_wysiwyg = "true";
defparam \xordvalue[8] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \xordvalue[1] (
	.clk(clk),
	.d(\xordvalue~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[1]~q ),
	.prn(vcc));
defparam \xordvalue[1] .is_wysiwyg = "true";
defparam \xordvalue[1] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \xordvalue[2] (
	.clk(clk),
	.d(\xordvalue~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[2]~q ),
	.prn(vcc));
defparam \xordvalue[2] .is_wysiwyg = "true";
defparam \xordvalue[2] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \xordvalue[3] (
	.clk(clk),
	.d(\xordvalue~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[3]~q ),
	.prn(vcc));
defparam \xordvalue[3] .is_wysiwyg = "true";
defparam \xordvalue[3] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \xordvalue[4] (
	.clk(clk),
	.d(\xordvalue~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[4]~q ),
	.prn(vcc));
defparam \xordvalue[4] .is_wysiwyg = "true";
defparam \xordvalue[4] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \xordvalue[5] (
	.clk(clk),
	.d(\xordvalue~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[5]~q ),
	.prn(vcc));
defparam \xordvalue[5] .is_wysiwyg = "true";
defparam \xordvalue[5] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \xordvalue[6] (
	.clk(clk),
	.d(\xordvalue~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[6]~q ),
	.prn(vcc));
defparam \xordvalue[6] .is_wysiwyg = "true";
defparam \xordvalue[6] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \xordvalue[7] (
	.clk(clk),
	.d(\xordvalue~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[7]~q ),
	.prn(vcc));
defparam \xordvalue[7] .is_wysiwyg = "true";
defparam \xordvalue[7] .power_up = "low";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe16),
	.datae(gnd),
	.dataf(!pipeline_dffe_01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~37 .shared_arith = "off";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h00000000000000FF;
defparam \Add0~41 .shared_arith = "off";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_18),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h00000000000000FF;
defparam \Add0~45 .shared_arith = "off";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout());
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h00000000000000FF;
defparam \Add0~49 .shared_arith = "off";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout());
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h00000000000000FF;
defparam \Add0~53 .shared_arith = "off";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout());
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h00000000000000FF;
defparam \Add0~57 .shared_arith = "off";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout());
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h00000000000000FF;
defparam \Add0~61 .shared_arith = "off";

arriav_lcell_comb \Add0~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~65_sumout ),
	.cout(\Add0~66 ),
	.shareout());
defparam \Add0~65 .extended_lut = "off";
defparam \Add0~65 .lut_mask = 64'h00000000000000FF;
defparam \Add0~65 .shared_arith = "off";

arriav_lcell_comb \Add0~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~69_sumout ),
	.cout(\Add0~70 ),
	.shareout());
defparam \Add0~69 .extended_lut = "off";
defparam \Add0~69 .lut_mask = 64'h00000000000000FF;
defparam \Add0~69 .shared_arith = "off";

arriav_lcell_comb \xordvalue~0 (
	.dataa(!dffe18),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

arriav_lcell_comb \xordvalue~1 (
	.dataa(!dffe9),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~1 .extended_lut = "off";
defparam \xordvalue~1 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~1 .shared_arith = "off";

arriav_lcell_comb \xordvalue~2 (
	.dataa(!dffe17),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~2 .extended_lut = "off";
defparam \xordvalue~2 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~2 .shared_arith = "off";

arriav_lcell_comb \xordvalue~3 (
	.dataa(!dffe10),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~3 .extended_lut = "off";
defparam \xordvalue~3 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~3 .shared_arith = "off";

arriav_lcell_comb \xordvalue~4 (
	.dataa(!dffe11),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~4 .extended_lut = "off";
defparam \xordvalue~4 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~4 .shared_arith = "off";

arriav_lcell_comb \xordvalue~5 (
	.dataa(!dffe12),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~5 .extended_lut = "off";
defparam \xordvalue~5 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~5 .shared_arith = "off";

arriav_lcell_comb \xordvalue~6 (
	.dataa(!dffe13),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~6 .extended_lut = "off";
defparam \xordvalue~6 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~6 .shared_arith = "off";

arriav_lcell_comb \xordvalue~7 (
	.dataa(!dffe14),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~7 .extended_lut = "off";
defparam \xordvalue~7 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~7 .shared_arith = "off";

arriav_lcell_comb \xordvalue~8 (
	.dataa(!dffe15),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~8 .extended_lut = "off";
defparam \xordvalue~8 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~8 .shared_arith = "off";

arriav_lcell_comb \xordvalue~9 (
	.dataa(!dffe161),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~9 .extended_lut = "off";
defparam \xordvalue~9 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~9 .shared_arith = "off";

endmodule

module nco_test_lpm_add_sub_7 (
	a_17,
	xordvalue_10,
	a_16,
	a_15,
	a_14,
	a_13,
	a_12,
	a_11,
	a_10,
	a_9,
	a_0,
	xordvalue_0,
	a_8,
	xordvalue_8,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	a_4,
	xordvalue_4,
	a_5,
	xordvalue_5,
	a_6,
	xordvalue_6,
	a_7,
	xordvalue_7,
	pipeline_dffe_17,
	pipeline_dffe_16,
	pipeline_dffe_15,
	pipeline_dffe_14,
	pipeline_dffe_13,
	pipeline_dffe_12,
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_9,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_10;
input 	a_16;
input 	a_15;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_10;
input 	a_9;
input 	a_0;
input 	xordvalue_0;
input 	a_8;
input 	xordvalue_8;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
input 	a_4;
input 	xordvalue_4;
input 	a_5;
input 	xordvalue_5;
input 	a_6;
input 	xordvalue_6;
input 	a_7;
input 	xordvalue_7;
output 	pipeline_dffe_17;
output 	pipeline_dffe_16;
output 	pipeline_dffe_15;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
output 	pipeline_dffe_9;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_add_sub_0qg_5 auto_generated(
	.a_17(a_17),
	.xordvalue_10(xordvalue_10),
	.a_16(a_16),
	.a_15(a_15),
	.a_14(a_14),
	.a_13(a_13),
	.a_12(a_12),
	.a_11(a_11),
	.a_10(a_10),
	.a_9(a_9),
	.a_0(a_0),
	.xordvalue_0(xordvalue_0),
	.a_8(a_8),
	.xordvalue_8(xordvalue_8),
	.a_1(a_1),
	.xordvalue_1(xordvalue_1),
	.a_2(a_2),
	.xordvalue_2(xordvalue_2),
	.a_3(a_3),
	.xordvalue_3(xordvalue_3),
	.a_4(a_4),
	.xordvalue_4(xordvalue_4),
	.a_5(a_5),
	.xordvalue_5(xordvalue_5),
	.a_6(a_6),
	.xordvalue_6(xordvalue_6),
	.a_7(a_7),
	.xordvalue_7(xordvalue_7),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module nco_test_add_sub_0qg_5 (
	a_17,
	xordvalue_10,
	a_16,
	a_15,
	a_14,
	a_13,
	a_12,
	a_11,
	a_10,
	a_9,
	a_0,
	xordvalue_0,
	a_8,
	xordvalue_8,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	a_4,
	xordvalue_4,
	a_5,
	xordvalue_5,
	a_6,
	xordvalue_6,
	a_7,
	xordvalue_7,
	pipeline_dffe_17,
	pipeline_dffe_16,
	pipeline_dffe_15,
	pipeline_dffe_14,
	pipeline_dffe_13,
	pipeline_dffe_12,
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_9,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_10;
input 	a_16;
input 	a_15;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_10;
input 	a_9;
input 	a_0;
input 	xordvalue_0;
input 	a_8;
input 	xordvalue_8;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
input 	a_4;
input 	xordvalue_4;
input 	a_5;
input 	xordvalue_5;
input 	a_6;
input 	xordvalue_6;
input 	a_7;
input 	xordvalue_7;
output 	pipeline_dffe_17;
output 	pipeline_dffe_16;
output 	pipeline_dffe_15;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
output 	pipeline_dffe_9;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \op_1~38 ;
wire \op_1~46 ;
wire \op_1~50 ;
wire \op_1~54 ;
wire \op_1~58 ;
wire \op_1~62 ;
wire \op_1~66 ;
wire \op_1~70 ;
wire \op_1~42 ;
wire \op_1~34 ;
wire \op_1~30 ;
wire \op_1~26 ;
wire \op_1~22 ;
wire \op_1~18 ;
wire \op_1~14 ;
wire \op_1~10 ;
wire \op_1~6 ;
wire \op_1~1_sumout ;
wire \op_1~5_sumout ;
wire \op_1~9_sumout ;
wire \op_1~13_sumout ;
wire \op_1~17_sumout ;
wire \op_1~21_sumout ;
wire \op_1~25_sumout ;
wire \op_1~29_sumout ;
wire \op_1~33_sumout ;
wire \op_1~37_sumout ;
wire \op_1~45_sumout ;
wire \op_1~49_sumout ;
wire \op_1~53_sumout ;
wire \op_1~57_sumout ;
wire \op_1~61_sumout ;
wire \op_1~65_sumout ;
wire \op_1~69_sumout ;
wire \op_1~41_sumout ;


dffeas \pipeline_dffe[17] (
	.clk(clock),
	.d(\op_1~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_17),
	.prn(vcc));
defparam \pipeline_dffe[17] .is_wysiwyg = "true";
defparam \pipeline_dffe[17] .power_up = "low";

dffeas \pipeline_dffe[16] (
	.clk(clock),
	.d(\op_1~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_16),
	.prn(vcc));
defparam \pipeline_dffe[16] .is_wysiwyg = "true";
defparam \pipeline_dffe[16] .power_up = "low";

dffeas \pipeline_dffe[15] (
	.clk(clock),
	.d(\op_1~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_15),
	.prn(vcc));
defparam \pipeline_dffe[15] .is_wysiwyg = "true";
defparam \pipeline_dffe[15] .power_up = "low";

dffeas \pipeline_dffe[14] (
	.clk(clock),
	.d(\op_1~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_14),
	.prn(vcc));
defparam \pipeline_dffe[14] .is_wysiwyg = "true";
defparam \pipeline_dffe[14] .power_up = "low";

dffeas \pipeline_dffe[13] (
	.clk(clock),
	.d(\op_1~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_13),
	.prn(vcc));
defparam \pipeline_dffe[13] .is_wysiwyg = "true";
defparam \pipeline_dffe[13] .power_up = "low";

dffeas \pipeline_dffe[12] (
	.clk(clock),
	.d(\op_1~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_12),
	.prn(vcc));
defparam \pipeline_dffe[12] .is_wysiwyg = "true";
defparam \pipeline_dffe[12] .power_up = "low";

dffeas \pipeline_dffe[11] (
	.clk(clock),
	.d(\op_1~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \pipeline_dffe[11] .is_wysiwyg = "true";
defparam \pipeline_dffe[11] .power_up = "low";

dffeas \pipeline_dffe[10] (
	.clk(clock),
	.d(\op_1~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \pipeline_dffe[10] .is_wysiwyg = "true";
defparam \pipeline_dffe[10] .power_up = "low";

dffeas \pipeline_dffe[9] (
	.clk(clock),
	.d(\op_1~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \pipeline_dffe[9] .is_wysiwyg = "true";
defparam \pipeline_dffe[9] .power_up = "low";

dffeas \pipeline_dffe[0] (
	.clk(clock),
	.d(\op_1~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_0),
	.prn(vcc));
defparam \pipeline_dffe[0] .is_wysiwyg = "true";
defparam \pipeline_dffe[0] .power_up = "low";

dffeas \pipeline_dffe[1] (
	.clk(clock),
	.d(\op_1~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_1),
	.prn(vcc));
defparam \pipeline_dffe[1] .is_wysiwyg = "true";
defparam \pipeline_dffe[1] .power_up = "low";

dffeas \pipeline_dffe[2] (
	.clk(clock),
	.d(\op_1~49_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \pipeline_dffe[2] .is_wysiwyg = "true";
defparam \pipeline_dffe[2] .power_up = "low";

dffeas \pipeline_dffe[3] (
	.clk(clock),
	.d(\op_1~53_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \pipeline_dffe[3] .is_wysiwyg = "true";
defparam \pipeline_dffe[3] .power_up = "low";

dffeas \pipeline_dffe[4] (
	.clk(clock),
	.d(\op_1~57_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \pipeline_dffe[4] .is_wysiwyg = "true";
defparam \pipeline_dffe[4] .power_up = "low";

dffeas \pipeline_dffe[5] (
	.clk(clock),
	.d(\op_1~61_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \pipeline_dffe[5] .is_wysiwyg = "true";
defparam \pipeline_dffe[5] .power_up = "low";

dffeas \pipeline_dffe[6] (
	.clk(clock),
	.d(\op_1~65_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \pipeline_dffe[6] .is_wysiwyg = "true";
defparam \pipeline_dffe[6] .power_up = "low";

dffeas \pipeline_dffe[7] (
	.clk(clock),
	.d(\op_1~69_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \pipeline_dffe[7] .is_wysiwyg = "true";
defparam \pipeline_dffe[7] .power_up = "low";

dffeas \pipeline_dffe[8] (
	.clk(clock),
	.d(\op_1~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \pipeline_dffe[8] .is_wysiwyg = "true";
defparam \pipeline_dffe[8] .power_up = "low";

arriav_lcell_comb \op_1~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~37_sumout ),
	.cout(\op_1~38 ),
	.shareout());
defparam \op_1~37 .extended_lut = "off";
defparam \op_1~37 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~37 .shared_arith = "off";

arriav_lcell_comb \op_1~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_1),
	.datag(gnd),
	.cin(\op_1~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~45_sumout ),
	.cout(\op_1~46 ),
	.shareout());
defparam \op_1~45 .extended_lut = "off";
defparam \op_1~45 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~45 .shared_arith = "off";

arriav_lcell_comb \op_1~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_2),
	.datag(gnd),
	.cin(\op_1~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~49_sumout ),
	.cout(\op_1~50 ),
	.shareout());
defparam \op_1~49 .extended_lut = "off";
defparam \op_1~49 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~49 .shared_arith = "off";

arriav_lcell_comb \op_1~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_3),
	.datag(gnd),
	.cin(\op_1~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~53_sumout ),
	.cout(\op_1~54 ),
	.shareout());
defparam \op_1~53 .extended_lut = "off";
defparam \op_1~53 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~53 .shared_arith = "off";

arriav_lcell_comb \op_1~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_4),
	.datag(gnd),
	.cin(\op_1~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~57_sumout ),
	.cout(\op_1~58 ),
	.shareout());
defparam \op_1~57 .extended_lut = "off";
defparam \op_1~57 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~57 .shared_arith = "off";

arriav_lcell_comb \op_1~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_5),
	.datag(gnd),
	.cin(\op_1~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~61_sumout ),
	.cout(\op_1~62 ),
	.shareout());
defparam \op_1~61 .extended_lut = "off";
defparam \op_1~61 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~61 .shared_arith = "off";

arriav_lcell_comb \op_1~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_6),
	.datag(gnd),
	.cin(\op_1~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~65_sumout ),
	.cout(\op_1~66 ),
	.shareout());
defparam \op_1~65 .extended_lut = "off";
defparam \op_1~65 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~65 .shared_arith = "off";

arriav_lcell_comb \op_1~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_7),
	.datag(gnd),
	.cin(\op_1~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~69_sumout ),
	.cout(\op_1~70 ),
	.shareout());
defparam \op_1~69 .extended_lut = "off";
defparam \op_1~69 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~69 .shared_arith = "off";

arriav_lcell_comb \op_1~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_8),
	.datag(gnd),
	.cin(\op_1~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~41_sumout ),
	.cout(\op_1~42 ),
	.shareout());
defparam \op_1~41 .extended_lut = "off";
defparam \op_1~41 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~41 .shared_arith = "off";

arriav_lcell_comb \op_1~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~33_sumout ),
	.cout(\op_1~34 ),
	.shareout());
defparam \op_1~33 .extended_lut = "off";
defparam \op_1~33 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~33 .shared_arith = "off";

arriav_lcell_comb \op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~29_sumout ),
	.cout(\op_1~30 ),
	.shareout());
defparam \op_1~29 .extended_lut = "off";
defparam \op_1~29 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~29 .shared_arith = "off";

arriav_lcell_comb \op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~25_sumout ),
	.cout(\op_1~26 ),
	.shareout());
defparam \op_1~25 .extended_lut = "off";
defparam \op_1~25 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~25 .shared_arith = "off";

arriav_lcell_comb \op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~21_sumout ),
	.cout(\op_1~22 ),
	.shareout());
defparam \op_1~21 .extended_lut = "off";
defparam \op_1~21 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~21 .shared_arith = "off";

arriav_lcell_comb \op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~17_sumout ),
	.cout(\op_1~18 ),
	.shareout());
defparam \op_1~17 .extended_lut = "off";
defparam \op_1~17 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~17 .shared_arith = "off";

arriav_lcell_comb \op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~13_sumout ),
	.cout(\op_1~14 ),
	.shareout());
defparam \op_1~13 .extended_lut = "off";
defparam \op_1~13 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~13 .shared_arith = "off";

arriav_lcell_comb \op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~9_sumout ),
	.cout(\op_1~10 ),
	.shareout());
defparam \op_1~9 .extended_lut = "off";
defparam \op_1~9 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~9 .shared_arith = "off";

arriav_lcell_comb \op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_16),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~5_sumout ),
	.cout(\op_1~6 ),
	.shareout());
defparam \op_1~5 .extended_lut = "off";
defparam \op_1~5 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~5 .shared_arith = "off";

arriav_lcell_comb \op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_17),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~1_sumout ),
	.cout(),
	.shareout());
defparam \op_1~1 .extended_lut = "off";
defparam \op_1~1 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~1 .shared_arith = "off";

endmodule

module nco_test_cordic_axor_1p_lpm_6 (
	sin_o_0,
	pipeline_dffe_17,
	pipeline_dffe_16,
	dffe16,
	dffe18,
	pipeline_dffe_15,
	pipeline_dffe_171,
	pipeline_dffe_14,
	pipeline_dffe_161,
	pipeline_dffe_13,
	dffe17,
	pipeline_dffe_151,
	pipeline_dffe_12,
	dffe161,
	pipeline_dffe_141,
	pipeline_dffe_10,
	pipeline_dffe_11,
	dffe15,
	pipeline_dffe_0,
	pipeline_dffe_131,
	dffe14,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_121,
	dffe13,
	pipeline_dffe_111,
	dffe12,
	dffe10,
	dffe11,
	pipeline_dffe_101,
	pipeline_dffe_91,
	pipeline_dffe_01,
	pipeline_dffe_18,
	pipeline_dffe_21,
	pipeline_dffe_31,
	pipeline_dffe_41,
	pipeline_dffe_51,
	pipeline_dffe_61,
	pipeline_dffe_71,
	pipeline_dffe_81,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	sin_o_0;
output 	pipeline_dffe_17;
output 	pipeline_dffe_16;
input 	dffe16;
input 	dffe18;
output 	pipeline_dffe_15;
input 	pipeline_dffe_171;
output 	pipeline_dffe_14;
input 	pipeline_dffe_161;
output 	pipeline_dffe_13;
input 	dffe17;
input 	pipeline_dffe_151;
output 	pipeline_dffe_12;
input 	dffe161;
input 	pipeline_dffe_141;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
input 	dffe15;
output 	pipeline_dffe_0;
input 	pipeline_dffe_131;
input 	dffe14;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	pipeline_dffe_121;
input 	dffe13;
input 	pipeline_dffe_111;
input 	dffe12;
input 	dffe10;
input 	dffe11;
input 	pipeline_dffe_101;
input 	pipeline_dffe_91;
input 	pipeline_dffe_01;
input 	pipeline_dffe_18;
input 	pipeline_dffe_21;
input 	pipeline_dffe_31;
input 	pipeline_dffe_41;
input 	pipeline_dffe_51;
input 	pipeline_dffe_61;
input 	pipeline_dffe_71;
input 	pipeline_dffe_81;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[17]~q ;
wire \xordvalue[10]~q ;
wire \Add0~1_sumout ;
wire \a[16]~q ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \a[15]~q ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \a[14]~q ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \a[13]~q ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \a[12]~q ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \a[11]~q ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \a[10]~q ;
wire \a[0]~q ;
wire \xordvalue[0]~q ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \a[9]~q ;
wire \a[1]~q ;
wire \xordvalue[1]~q ;
wire \a[2]~q ;
wire \xordvalue[2]~q ;
wire \a[3]~q ;
wire \xordvalue[3]~q ;
wire \a[4]~q ;
wire \xordvalue[4]~q ;
wire \a[5]~q ;
wire \xordvalue[5]~q ;
wire \a[6]~q ;
wire \xordvalue[6]~q ;
wire \a[7]~q ;
wire \xordvalue[7]~q ;
wire \a[8]~q ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~65_sumout ;
wire \Add0~66 ;
wire \Add0~69_sumout ;
wire \Add0~70 ;
wire \xordvalue~0_combout ;
wire \xordvalue~1_combout ;
wire \xordvalue~2_combout ;
wire \xordvalue~3_combout ;
wire \xordvalue~4_combout ;
wire \xordvalue~5_combout ;
wire \xordvalue~6_combout ;
wire \xordvalue~7_combout ;
wire \xordvalue~8_combout ;


nco_test_lpm_add_sub_8 u0(
	.a_17(\a[17]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.a_16(\a[16]~q ),
	.a_15(\a[15]~q ),
	.a_14(\a[14]~q ),
	.a_13(\a[13]~q ),
	.a_12(\a[12]~q ),
	.a_11(\a[11]~q ),
	.a_10(\a[10]~q ),
	.a_0(\a[0]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_9(\a[9]~q ),
	.a_1(\a[1]~q ),
	.xordvalue_1(\xordvalue[1]~q ),
	.a_2(\a[2]~q ),
	.xordvalue_2(\xordvalue[2]~q ),
	.a_3(\a[3]~q ),
	.xordvalue_3(\xordvalue[3]~q ),
	.a_4(\a[4]~q ),
	.xordvalue_4(\xordvalue[4]~q ),
	.a_5(\a[5]~q ),
	.xordvalue_5(\xordvalue[5]~q ),
	.a_6(\a[6]~q ),
	.xordvalue_6(\xordvalue[6]~q ),
	.a_7(\a[7]~q ),
	.xordvalue_7(\xordvalue[7]~q ),
	.a_8(\a[8]~q ),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[17] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[17]~q ),
	.prn(vcc));
defparam \a[17] .is_wysiwyg = "true";
defparam \a[17] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_171),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h00000000000000FF;
defparam \Add0~1 .shared_arith = "off";

dffeas \a[16] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[16]~q ),
	.prn(vcc));
defparam \a[16] .is_wysiwyg = "true";
defparam \a[16] .power_up = "low";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h00000000000000FF;
defparam \Add0~5 .shared_arith = "off";

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h00000000000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h00000000000000FF;
defparam \Add0~13 .shared_arith = "off";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h00000000000000FF;
defparam \Add0~17 .shared_arith = "off";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h00000000000000FF;
defparam \Add0~21 .shared_arith = "off";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h00000000000000FF;
defparam \Add0~25 .shared_arith = "off";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h00000000000000FF;
defparam \Add0~29 .shared_arith = "off";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \xordvalue[1] (
	.clk(clk),
	.d(\xordvalue~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[1]~q ),
	.prn(vcc));
defparam \xordvalue[1] .is_wysiwyg = "true";
defparam \xordvalue[1] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \xordvalue[2] (
	.clk(clk),
	.d(\xordvalue~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[2]~q ),
	.prn(vcc));
defparam \xordvalue[2] .is_wysiwyg = "true";
defparam \xordvalue[2] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \xordvalue[3] (
	.clk(clk),
	.d(\xordvalue~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[3]~q ),
	.prn(vcc));
defparam \xordvalue[3] .is_wysiwyg = "true";
defparam \xordvalue[3] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \xordvalue[4] (
	.clk(clk),
	.d(\xordvalue~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[4]~q ),
	.prn(vcc));
defparam \xordvalue[4] .is_wysiwyg = "true";
defparam \xordvalue[4] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \xordvalue[5] (
	.clk(clk),
	.d(\xordvalue~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[5]~q ),
	.prn(vcc));
defparam \xordvalue[5] .is_wysiwyg = "true";
defparam \xordvalue[5] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \xordvalue[6] (
	.clk(clk),
	.d(\xordvalue~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[6]~q ),
	.prn(vcc));
defparam \xordvalue[6] .is_wysiwyg = "true";
defparam \xordvalue[6] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \xordvalue[7] (
	.clk(clk),
	.d(\xordvalue~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[7]~q ),
	.prn(vcc));
defparam \xordvalue[7] .is_wysiwyg = "true";
defparam \xordvalue[7] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe16),
	.datae(gnd),
	.dataf(!pipeline_dffe_01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~33 .shared_arith = "off";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h00000000000000FF;
defparam \Add0~37 .shared_arith = "off";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_18),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h00000000000000FF;
defparam \Add0~41 .shared_arith = "off";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h00000000000000FF;
defparam \Add0~45 .shared_arith = "off";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout());
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h00000000000000FF;
defparam \Add0~49 .shared_arith = "off";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout());
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h00000000000000FF;
defparam \Add0~53 .shared_arith = "off";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout());
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h00000000000000FF;
defparam \Add0~57 .shared_arith = "off";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout());
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h00000000000000FF;
defparam \Add0~61 .shared_arith = "off";

arriav_lcell_comb \Add0~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~65_sumout ),
	.cout(\Add0~66 ),
	.shareout());
defparam \Add0~65 .extended_lut = "off";
defparam \Add0~65 .lut_mask = 64'h00000000000000FF;
defparam \Add0~65 .shared_arith = "off";

arriav_lcell_comb \Add0~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~69_sumout ),
	.cout(\Add0~70 ),
	.shareout());
defparam \Add0~69 .extended_lut = "off";
defparam \Add0~69 .lut_mask = 64'h00000000000000FF;
defparam \Add0~69 .shared_arith = "off";

arriav_lcell_comb \xordvalue~0 (
	.dataa(!dffe16),
	.datab(!dffe18),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

arriav_lcell_comb \xordvalue~1 (
	.dataa(!dffe16),
	.datab(!dffe10),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~1 .extended_lut = "off";
defparam \xordvalue~1 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~1 .shared_arith = "off";

arriav_lcell_comb \xordvalue~2 (
	.dataa(!dffe16),
	.datab(!dffe11),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~2 .extended_lut = "off";
defparam \xordvalue~2 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~2 .shared_arith = "off";

arriav_lcell_comb \xordvalue~3 (
	.dataa(!dffe16),
	.datab(!dffe12),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~3 .extended_lut = "off";
defparam \xordvalue~3 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~3 .shared_arith = "off";

arriav_lcell_comb \xordvalue~4 (
	.dataa(!dffe16),
	.datab(!dffe13),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~4 .extended_lut = "off";
defparam \xordvalue~4 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~4 .shared_arith = "off";

arriav_lcell_comb \xordvalue~5 (
	.dataa(!dffe16),
	.datab(!dffe14),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~5 .extended_lut = "off";
defparam \xordvalue~5 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~5 .shared_arith = "off";

arriav_lcell_comb \xordvalue~6 (
	.dataa(!dffe16),
	.datab(!dffe15),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~6 .extended_lut = "off";
defparam \xordvalue~6 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~6 .shared_arith = "off";

arriav_lcell_comb \xordvalue~7 (
	.dataa(!dffe16),
	.datab(!dffe161),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~7 .extended_lut = "off";
defparam \xordvalue~7 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~7 .shared_arith = "off";

arriav_lcell_comb \xordvalue~8 (
	.dataa(!dffe16),
	.datab(!dffe17),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~8 .extended_lut = "off";
defparam \xordvalue~8 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~8 .shared_arith = "off";

endmodule

module nco_test_lpm_add_sub_8 (
	a_17,
	xordvalue_10,
	a_16,
	a_15,
	a_14,
	a_13,
	a_12,
	a_11,
	a_10,
	a_0,
	xordvalue_0,
	a_9,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	a_4,
	xordvalue_4,
	a_5,
	xordvalue_5,
	a_6,
	xordvalue_6,
	a_7,
	xordvalue_7,
	a_8,
	pipeline_dffe_17,
	pipeline_dffe_16,
	pipeline_dffe_15,
	pipeline_dffe_14,
	pipeline_dffe_13,
	pipeline_dffe_12,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_10;
input 	a_16;
input 	a_15;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_10;
input 	a_0;
input 	xordvalue_0;
input 	a_9;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
input 	a_4;
input 	xordvalue_4;
input 	a_5;
input 	xordvalue_5;
input 	a_6;
input 	xordvalue_6;
input 	a_7;
input 	xordvalue_7;
input 	a_8;
output 	pipeline_dffe_17;
output 	pipeline_dffe_16;
output 	pipeline_dffe_15;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
output 	pipeline_dffe_12;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_add_sub_0qg_6 auto_generated(
	.a_17(a_17),
	.xordvalue_10(xordvalue_10),
	.a_16(a_16),
	.a_15(a_15),
	.a_14(a_14),
	.a_13(a_13),
	.a_12(a_12),
	.a_11(a_11),
	.a_10(a_10),
	.a_0(a_0),
	.xordvalue_0(xordvalue_0),
	.a_9(a_9),
	.a_1(a_1),
	.xordvalue_1(xordvalue_1),
	.a_2(a_2),
	.xordvalue_2(xordvalue_2),
	.a_3(a_3),
	.xordvalue_3(xordvalue_3),
	.a_4(a_4),
	.xordvalue_4(xordvalue_4),
	.a_5(a_5),
	.xordvalue_5(xordvalue_5),
	.a_6(a_6),
	.xordvalue_6(xordvalue_6),
	.a_7(a_7),
	.xordvalue_7(xordvalue_7),
	.a_8(a_8),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module nco_test_add_sub_0qg_6 (
	a_17,
	xordvalue_10,
	a_16,
	a_15,
	a_14,
	a_13,
	a_12,
	a_11,
	a_10,
	a_0,
	xordvalue_0,
	a_9,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	a_4,
	xordvalue_4,
	a_5,
	xordvalue_5,
	a_6,
	xordvalue_6,
	a_7,
	xordvalue_7,
	a_8,
	pipeline_dffe_17,
	pipeline_dffe_16,
	pipeline_dffe_15,
	pipeline_dffe_14,
	pipeline_dffe_13,
	pipeline_dffe_12,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_10;
input 	a_16;
input 	a_15;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_10;
input 	a_0;
input 	xordvalue_0;
input 	a_9;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
input 	a_4;
input 	xordvalue_4;
input 	a_5;
input 	xordvalue_5;
input 	a_6;
input 	xordvalue_6;
input 	a_7;
input 	xordvalue_7;
input 	a_8;
output 	pipeline_dffe_17;
output 	pipeline_dffe_16;
output 	pipeline_dffe_15;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
output 	pipeline_dffe_12;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \op_1~34 ;
wire \op_1~42 ;
wire \op_1~46 ;
wire \op_1~50 ;
wire \op_1~54 ;
wire \op_1~58 ;
wire \op_1~62 ;
wire \op_1~66 ;
wire \op_1~70 ;
wire \op_1~38 ;
wire \op_1~30 ;
wire \op_1~26 ;
wire \op_1~22 ;
wire \op_1~18 ;
wire \op_1~14 ;
wire \op_1~10 ;
wire \op_1~6 ;
wire \op_1~1_sumout ;
wire \op_1~5_sumout ;
wire \op_1~9_sumout ;
wire \op_1~13_sumout ;
wire \op_1~17_sumout ;
wire \op_1~21_sumout ;
wire \op_1~29_sumout ;
wire \op_1~25_sumout ;
wire \op_1~33_sumout ;
wire \op_1~41_sumout ;
wire \op_1~45_sumout ;
wire \op_1~49_sumout ;
wire \op_1~53_sumout ;
wire \op_1~57_sumout ;
wire \op_1~61_sumout ;
wire \op_1~65_sumout ;
wire \op_1~69_sumout ;
wire \op_1~37_sumout ;


dffeas \pipeline_dffe[17] (
	.clk(clock),
	.d(\op_1~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_17),
	.prn(vcc));
defparam \pipeline_dffe[17] .is_wysiwyg = "true";
defparam \pipeline_dffe[17] .power_up = "low";

dffeas \pipeline_dffe[16] (
	.clk(clock),
	.d(\op_1~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_16),
	.prn(vcc));
defparam \pipeline_dffe[16] .is_wysiwyg = "true";
defparam \pipeline_dffe[16] .power_up = "low";

dffeas \pipeline_dffe[15] (
	.clk(clock),
	.d(\op_1~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_15),
	.prn(vcc));
defparam \pipeline_dffe[15] .is_wysiwyg = "true";
defparam \pipeline_dffe[15] .power_up = "low";

dffeas \pipeline_dffe[14] (
	.clk(clock),
	.d(\op_1~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_14),
	.prn(vcc));
defparam \pipeline_dffe[14] .is_wysiwyg = "true";
defparam \pipeline_dffe[14] .power_up = "low";

dffeas \pipeline_dffe[13] (
	.clk(clock),
	.d(\op_1~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_13),
	.prn(vcc));
defparam \pipeline_dffe[13] .is_wysiwyg = "true";
defparam \pipeline_dffe[13] .power_up = "low";

dffeas \pipeline_dffe[12] (
	.clk(clock),
	.d(\op_1~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_12),
	.prn(vcc));
defparam \pipeline_dffe[12] .is_wysiwyg = "true";
defparam \pipeline_dffe[12] .power_up = "low";

dffeas \pipeline_dffe[10] (
	.clk(clock),
	.d(\op_1~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \pipeline_dffe[10] .is_wysiwyg = "true";
defparam \pipeline_dffe[10] .power_up = "low";

dffeas \pipeline_dffe[11] (
	.clk(clock),
	.d(\op_1~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \pipeline_dffe[11] .is_wysiwyg = "true";
defparam \pipeline_dffe[11] .power_up = "low";

dffeas \pipeline_dffe[0] (
	.clk(clock),
	.d(\op_1~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_0),
	.prn(vcc));
defparam \pipeline_dffe[0] .is_wysiwyg = "true";
defparam \pipeline_dffe[0] .power_up = "low";

dffeas \pipeline_dffe[1] (
	.clk(clock),
	.d(\op_1~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_1),
	.prn(vcc));
defparam \pipeline_dffe[1] .is_wysiwyg = "true";
defparam \pipeline_dffe[1] .power_up = "low";

dffeas \pipeline_dffe[2] (
	.clk(clock),
	.d(\op_1~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \pipeline_dffe[2] .is_wysiwyg = "true";
defparam \pipeline_dffe[2] .power_up = "low";

dffeas \pipeline_dffe[3] (
	.clk(clock),
	.d(\op_1~49_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \pipeline_dffe[3] .is_wysiwyg = "true";
defparam \pipeline_dffe[3] .power_up = "low";

dffeas \pipeline_dffe[4] (
	.clk(clock),
	.d(\op_1~53_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \pipeline_dffe[4] .is_wysiwyg = "true";
defparam \pipeline_dffe[4] .power_up = "low";

dffeas \pipeline_dffe[5] (
	.clk(clock),
	.d(\op_1~57_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \pipeline_dffe[5] .is_wysiwyg = "true";
defparam \pipeline_dffe[5] .power_up = "low";

dffeas \pipeline_dffe[6] (
	.clk(clock),
	.d(\op_1~61_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \pipeline_dffe[6] .is_wysiwyg = "true";
defparam \pipeline_dffe[6] .power_up = "low";

dffeas \pipeline_dffe[7] (
	.clk(clock),
	.d(\op_1~65_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \pipeline_dffe[7] .is_wysiwyg = "true";
defparam \pipeline_dffe[7] .power_up = "low";

dffeas \pipeline_dffe[8] (
	.clk(clock),
	.d(\op_1~69_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \pipeline_dffe[8] .is_wysiwyg = "true";
defparam \pipeline_dffe[8] .power_up = "low";

dffeas \pipeline_dffe[9] (
	.clk(clock),
	.d(\op_1~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \pipeline_dffe[9] .is_wysiwyg = "true";
defparam \pipeline_dffe[9] .power_up = "low";

arriav_lcell_comb \op_1~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~33_sumout ),
	.cout(\op_1~34 ),
	.shareout());
defparam \op_1~33 .extended_lut = "off";
defparam \op_1~33 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~33 .shared_arith = "off";

arriav_lcell_comb \op_1~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_1),
	.datag(gnd),
	.cin(\op_1~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~41_sumout ),
	.cout(\op_1~42 ),
	.shareout());
defparam \op_1~41 .extended_lut = "off";
defparam \op_1~41 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~41 .shared_arith = "off";

arriav_lcell_comb \op_1~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_2),
	.datag(gnd),
	.cin(\op_1~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~45_sumout ),
	.cout(\op_1~46 ),
	.shareout());
defparam \op_1~45 .extended_lut = "off";
defparam \op_1~45 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~45 .shared_arith = "off";

arriav_lcell_comb \op_1~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_3),
	.datag(gnd),
	.cin(\op_1~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~49_sumout ),
	.cout(\op_1~50 ),
	.shareout());
defparam \op_1~49 .extended_lut = "off";
defparam \op_1~49 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~49 .shared_arith = "off";

arriav_lcell_comb \op_1~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_4),
	.datag(gnd),
	.cin(\op_1~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~53_sumout ),
	.cout(\op_1~54 ),
	.shareout());
defparam \op_1~53 .extended_lut = "off";
defparam \op_1~53 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~53 .shared_arith = "off";

arriav_lcell_comb \op_1~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_5),
	.datag(gnd),
	.cin(\op_1~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~57_sumout ),
	.cout(\op_1~58 ),
	.shareout());
defparam \op_1~57 .extended_lut = "off";
defparam \op_1~57 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~57 .shared_arith = "off";

arriav_lcell_comb \op_1~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_6),
	.datag(gnd),
	.cin(\op_1~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~61_sumout ),
	.cout(\op_1~62 ),
	.shareout());
defparam \op_1~61 .extended_lut = "off";
defparam \op_1~61 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~61 .shared_arith = "off";

arriav_lcell_comb \op_1~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_7),
	.datag(gnd),
	.cin(\op_1~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~65_sumout ),
	.cout(\op_1~66 ),
	.shareout());
defparam \op_1~65 .extended_lut = "off";
defparam \op_1~65 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~65 .shared_arith = "off";

arriav_lcell_comb \op_1~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~69_sumout ),
	.cout(\op_1~70 ),
	.shareout());
defparam \op_1~69 .extended_lut = "off";
defparam \op_1~69 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~69 .shared_arith = "off";

arriav_lcell_comb \op_1~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~37_sumout ),
	.cout(\op_1~38 ),
	.shareout());
defparam \op_1~37 .extended_lut = "off";
defparam \op_1~37 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~37 .shared_arith = "off";

arriav_lcell_comb \op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~29_sumout ),
	.cout(\op_1~30 ),
	.shareout());
defparam \op_1~29 .extended_lut = "off";
defparam \op_1~29 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~29 .shared_arith = "off";

arriav_lcell_comb \op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~25_sumout ),
	.cout(\op_1~26 ),
	.shareout());
defparam \op_1~25 .extended_lut = "off";
defparam \op_1~25 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~25 .shared_arith = "off";

arriav_lcell_comb \op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~21_sumout ),
	.cout(\op_1~22 ),
	.shareout());
defparam \op_1~21 .extended_lut = "off";
defparam \op_1~21 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~21 .shared_arith = "off";

arriav_lcell_comb \op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~17_sumout ),
	.cout(\op_1~18 ),
	.shareout());
defparam \op_1~17 .extended_lut = "off";
defparam \op_1~17 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~17 .shared_arith = "off";

arriav_lcell_comb \op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~13_sumout ),
	.cout(\op_1~14 ),
	.shareout());
defparam \op_1~13 .extended_lut = "off";
defparam \op_1~13 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~13 .shared_arith = "off";

arriav_lcell_comb \op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~9_sumout ),
	.cout(\op_1~10 ),
	.shareout());
defparam \op_1~9 .extended_lut = "off";
defparam \op_1~9 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~9 .shared_arith = "off";

arriav_lcell_comb \op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_16),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~5_sumout ),
	.cout(\op_1~6 ),
	.shareout());
defparam \op_1~5 .extended_lut = "off";
defparam \op_1~5 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~5 .shared_arith = "off";

arriav_lcell_comb \op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_17),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~1_sumout ),
	.cout(),
	.shareout());
defparam \op_1~1 .extended_lut = "off";
defparam \op_1~1 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~1 .shared_arith = "off";

endmodule

module nco_test_cordic_axor_1p_lpm_7 (
	sin_o_0,
	pipeline_dffe_17,
	pipeline_dffe_16,
	dffe16,
	pipeline_dffe_15,
	pipeline_dffe_171,
	dffe18,
	pipeline_dffe_14,
	pipeline_dffe_13,
	dffe17,
	pipeline_dffe_161,
	pipeline_dffe_12,
	dffe161,
	pipeline_dffe_11,
	pipeline_dffe_151,
	pipeline_dffe_0,
	dffe15,
	pipeline_dffe_141,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	dffe14,
	pipeline_dffe_131,
	dffe13,
	pipeline_dffe_121,
	dffe11,
	dffe12,
	pipeline_dffe_101,
	pipeline_dffe_111,
	pipeline_dffe_01,
	pipeline_dffe_18,
	pipeline_dffe_21,
	pipeline_dffe_31,
	pipeline_dffe_41,
	pipeline_dffe_51,
	pipeline_dffe_61,
	pipeline_dffe_71,
	pipeline_dffe_81,
	pipeline_dffe_91,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	sin_o_0;
output 	pipeline_dffe_17;
output 	pipeline_dffe_16;
input 	dffe16;
output 	pipeline_dffe_15;
input 	pipeline_dffe_171;
input 	dffe18;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
input 	dffe17;
input 	pipeline_dffe_161;
output 	pipeline_dffe_12;
input 	dffe161;
output 	pipeline_dffe_11;
input 	pipeline_dffe_151;
output 	pipeline_dffe_0;
input 	dffe15;
input 	pipeline_dffe_141;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
input 	dffe14;
input 	pipeline_dffe_131;
input 	dffe13;
input 	pipeline_dffe_121;
input 	dffe11;
input 	dffe12;
input 	pipeline_dffe_101;
input 	pipeline_dffe_111;
input 	pipeline_dffe_01;
input 	pipeline_dffe_18;
input 	pipeline_dffe_21;
input 	pipeline_dffe_31;
input 	pipeline_dffe_41;
input 	pipeline_dffe_51;
input 	pipeline_dffe_61;
input 	pipeline_dffe_71;
input 	pipeline_dffe_81;
input 	pipeline_dffe_91;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[17]~q ;
wire \xordvalue[10]~q ;
wire \Add0~1_sumout ;
wire \a[16]~q ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \a[15]~q ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \a[14]~q ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \a[13]~q ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \a[12]~q ;
wire \a[11]~q ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \a[0]~q ;
wire \xordvalue[0]~q ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \a[10]~q ;
wire \a[1]~q ;
wire \xordvalue[1]~q ;
wire \a[2]~q ;
wire \xordvalue[2]~q ;
wire \a[3]~q ;
wire \xordvalue[3]~q ;
wire \a[4]~q ;
wire \xordvalue[4]~q ;
wire \a[5]~q ;
wire \xordvalue[5]~q ;
wire \a[6]~q ;
wire \xordvalue[6]~q ;
wire \a[7]~q ;
wire \a[8]~q ;
wire \a[9]~q ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~65_sumout ;
wire \Add0~66 ;
wire \Add0~69_sumout ;
wire \Add0~70 ;
wire \xordvalue~0_combout ;
wire \xordvalue~1_combout ;
wire \xordvalue~2_combout ;
wire \xordvalue~3_combout ;
wire \xordvalue~4_combout ;
wire \xordvalue~5_combout ;
wire \xordvalue~6_combout ;
wire \xordvalue~7_combout ;


nco_test_lpm_add_sub_9 u0(
	.a_17(\a[17]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.a_16(\a[16]~q ),
	.a_15(\a[15]~q ),
	.a_14(\a[14]~q ),
	.a_13(\a[13]~q ),
	.a_12(\a[12]~q ),
	.a_11(\a[11]~q ),
	.a_0(\a[0]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_10(\a[10]~q ),
	.a_1(\a[1]~q ),
	.xordvalue_1(\xordvalue[1]~q ),
	.a_2(\a[2]~q ),
	.xordvalue_2(\xordvalue[2]~q ),
	.a_3(\a[3]~q ),
	.xordvalue_3(\xordvalue[3]~q ),
	.a_4(\a[4]~q ),
	.xordvalue_4(\xordvalue[4]~q ),
	.a_5(\a[5]~q ),
	.xordvalue_5(\xordvalue[5]~q ),
	.a_6(\a[6]~q ),
	.xordvalue_6(\xordvalue[6]~q ),
	.a_7(\a[7]~q ),
	.a_8(\a[8]~q ),
	.a_9(\a[9]~q ),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[17] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[17]~q ),
	.prn(vcc));
defparam \a[17] .is_wysiwyg = "true";
defparam \a[17] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_171),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h00000000000000FF;
defparam \Add0~1 .shared_arith = "off";

dffeas \a[16] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[16]~q ),
	.prn(vcc));
defparam \a[16] .is_wysiwyg = "true";
defparam \a[16] .power_up = "low";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h00000000000000FF;
defparam \Add0~5 .shared_arith = "off";

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h00000000000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h00000000000000FF;
defparam \Add0~13 .shared_arith = "off";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h00000000000000FF;
defparam \Add0~17 .shared_arith = "off";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h00000000000000FF;
defparam \Add0~21 .shared_arith = "off";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h00000000000000FF;
defparam \Add0~25 .shared_arith = "off";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \xordvalue[1] (
	.clk(clk),
	.d(\xordvalue~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[1]~q ),
	.prn(vcc));
defparam \xordvalue[1] .is_wysiwyg = "true";
defparam \xordvalue[1] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \xordvalue[2] (
	.clk(clk),
	.d(\xordvalue~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[2]~q ),
	.prn(vcc));
defparam \xordvalue[2] .is_wysiwyg = "true";
defparam \xordvalue[2] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \xordvalue[3] (
	.clk(clk),
	.d(\xordvalue~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[3]~q ),
	.prn(vcc));
defparam \xordvalue[3] .is_wysiwyg = "true";
defparam \xordvalue[3] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \xordvalue[4] (
	.clk(clk),
	.d(\xordvalue~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[4]~q ),
	.prn(vcc));
defparam \xordvalue[4] .is_wysiwyg = "true";
defparam \xordvalue[4] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \xordvalue[5] (
	.clk(clk),
	.d(\xordvalue~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[5]~q ),
	.prn(vcc));
defparam \xordvalue[5] .is_wysiwyg = "true";
defparam \xordvalue[5] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \xordvalue[6] (
	.clk(clk),
	.d(\xordvalue~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[6]~q ),
	.prn(vcc));
defparam \xordvalue[6] .is_wysiwyg = "true";
defparam \xordvalue[6] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe16),
	.datae(gnd),
	.dataf(!pipeline_dffe_01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~29 .shared_arith = "off";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h00000000000000FF;
defparam \Add0~33 .shared_arith = "off";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_18),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h00000000000000FF;
defparam \Add0~37 .shared_arith = "off";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h00000000000000FF;
defparam \Add0~41 .shared_arith = "off";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h00000000000000FF;
defparam \Add0~45 .shared_arith = "off";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout());
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h00000000000000FF;
defparam \Add0~49 .shared_arith = "off";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout());
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h00000000000000FF;
defparam \Add0~53 .shared_arith = "off";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout());
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h00000000000000FF;
defparam \Add0~57 .shared_arith = "off";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout());
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h00000000000000FF;
defparam \Add0~61 .shared_arith = "off";

arriav_lcell_comb \Add0~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~65_sumout ),
	.cout(\Add0~66 ),
	.shareout());
defparam \Add0~65 .extended_lut = "off";
defparam \Add0~65 .lut_mask = 64'h00000000000000FF;
defparam \Add0~65 .shared_arith = "off";

arriav_lcell_comb \Add0~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~69_sumout ),
	.cout(\Add0~70 ),
	.shareout());
defparam \Add0~69 .extended_lut = "off";
defparam \Add0~69 .lut_mask = 64'h00000000000000FF;
defparam \Add0~69 .shared_arith = "off";

arriav_lcell_comb \xordvalue~0 (
	.dataa(!dffe18),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

arriav_lcell_comb \xordvalue~1 (
	.dataa(!dffe11),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~1 .extended_lut = "off";
defparam \xordvalue~1 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~1 .shared_arith = "off";

arriav_lcell_comb \xordvalue~2 (
	.dataa(!dffe12),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~2 .extended_lut = "off";
defparam \xordvalue~2 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~2 .shared_arith = "off";

arriav_lcell_comb \xordvalue~3 (
	.dataa(!dffe13),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~3 .extended_lut = "off";
defparam \xordvalue~3 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~3 .shared_arith = "off";

arriav_lcell_comb \xordvalue~4 (
	.dataa(!dffe14),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~4 .extended_lut = "off";
defparam \xordvalue~4 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~4 .shared_arith = "off";

arriav_lcell_comb \xordvalue~5 (
	.dataa(!dffe15),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~5 .extended_lut = "off";
defparam \xordvalue~5 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~5 .shared_arith = "off";

arriav_lcell_comb \xordvalue~6 (
	.dataa(!dffe161),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~6 .extended_lut = "off";
defparam \xordvalue~6 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~6 .shared_arith = "off";

arriav_lcell_comb \xordvalue~7 (
	.dataa(!dffe17),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~7 .extended_lut = "off";
defparam \xordvalue~7 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~7 .shared_arith = "off";

endmodule

module nco_test_lpm_add_sub_9 (
	a_17,
	xordvalue_10,
	a_16,
	a_15,
	a_14,
	a_13,
	a_12,
	a_11,
	a_0,
	xordvalue_0,
	a_10,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	a_4,
	xordvalue_4,
	a_5,
	xordvalue_5,
	a_6,
	xordvalue_6,
	a_7,
	a_8,
	a_9,
	pipeline_dffe_17,
	pipeline_dffe_16,
	pipeline_dffe_15,
	pipeline_dffe_14,
	pipeline_dffe_13,
	pipeline_dffe_12,
	pipeline_dffe_11,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_10;
input 	a_16;
input 	a_15;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_0;
input 	xordvalue_0;
input 	a_10;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
input 	a_4;
input 	xordvalue_4;
input 	a_5;
input 	xordvalue_5;
input 	a_6;
input 	xordvalue_6;
input 	a_7;
input 	a_8;
input 	a_9;
output 	pipeline_dffe_17;
output 	pipeline_dffe_16;
output 	pipeline_dffe_15;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_add_sub_0qg_7 auto_generated(
	.a_17(a_17),
	.xordvalue_10(xordvalue_10),
	.a_16(a_16),
	.a_15(a_15),
	.a_14(a_14),
	.a_13(a_13),
	.a_12(a_12),
	.a_11(a_11),
	.a_0(a_0),
	.xordvalue_0(xordvalue_0),
	.a_10(a_10),
	.a_1(a_1),
	.xordvalue_1(xordvalue_1),
	.a_2(a_2),
	.xordvalue_2(xordvalue_2),
	.a_3(a_3),
	.xordvalue_3(xordvalue_3),
	.a_4(a_4),
	.xordvalue_4(xordvalue_4),
	.a_5(a_5),
	.xordvalue_5(xordvalue_5),
	.a_6(a_6),
	.xordvalue_6(xordvalue_6),
	.a_7(a_7),
	.a_8(a_8),
	.a_9(a_9),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module nco_test_add_sub_0qg_7 (
	a_17,
	xordvalue_10,
	a_16,
	a_15,
	a_14,
	a_13,
	a_12,
	a_11,
	a_0,
	xordvalue_0,
	a_10,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	a_4,
	xordvalue_4,
	a_5,
	xordvalue_5,
	a_6,
	xordvalue_6,
	a_7,
	a_8,
	a_9,
	pipeline_dffe_17,
	pipeline_dffe_16,
	pipeline_dffe_15,
	pipeline_dffe_14,
	pipeline_dffe_13,
	pipeline_dffe_12,
	pipeline_dffe_11,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_10;
input 	a_16;
input 	a_15;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_0;
input 	xordvalue_0;
input 	a_10;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
input 	a_4;
input 	xordvalue_4;
input 	a_5;
input 	xordvalue_5;
input 	a_6;
input 	xordvalue_6;
input 	a_7;
input 	a_8;
input 	a_9;
output 	pipeline_dffe_17;
output 	pipeline_dffe_16;
output 	pipeline_dffe_15;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \op_1~30 ;
wire \op_1~38 ;
wire \op_1~42 ;
wire \op_1~46 ;
wire \op_1~50 ;
wire \op_1~54 ;
wire \op_1~58 ;
wire \op_1~62 ;
wire \op_1~66 ;
wire \op_1~70 ;
wire \op_1~34 ;
wire \op_1~26 ;
wire \op_1~22 ;
wire \op_1~18 ;
wire \op_1~14 ;
wire \op_1~10 ;
wire \op_1~6 ;
wire \op_1~1_sumout ;
wire \op_1~5_sumout ;
wire \op_1~9_sumout ;
wire \op_1~13_sumout ;
wire \op_1~17_sumout ;
wire \op_1~21_sumout ;
wire \op_1~25_sumout ;
wire \op_1~29_sumout ;
wire \op_1~37_sumout ;
wire \op_1~41_sumout ;
wire \op_1~45_sumout ;
wire \op_1~49_sumout ;
wire \op_1~53_sumout ;
wire \op_1~57_sumout ;
wire \op_1~61_sumout ;
wire \op_1~65_sumout ;
wire \op_1~69_sumout ;
wire \op_1~33_sumout ;


dffeas \pipeline_dffe[17] (
	.clk(clock),
	.d(\op_1~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_17),
	.prn(vcc));
defparam \pipeline_dffe[17] .is_wysiwyg = "true";
defparam \pipeline_dffe[17] .power_up = "low";

dffeas \pipeline_dffe[16] (
	.clk(clock),
	.d(\op_1~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_16),
	.prn(vcc));
defparam \pipeline_dffe[16] .is_wysiwyg = "true";
defparam \pipeline_dffe[16] .power_up = "low";

dffeas \pipeline_dffe[15] (
	.clk(clock),
	.d(\op_1~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_15),
	.prn(vcc));
defparam \pipeline_dffe[15] .is_wysiwyg = "true";
defparam \pipeline_dffe[15] .power_up = "low";

dffeas \pipeline_dffe[14] (
	.clk(clock),
	.d(\op_1~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_14),
	.prn(vcc));
defparam \pipeline_dffe[14] .is_wysiwyg = "true";
defparam \pipeline_dffe[14] .power_up = "low";

dffeas \pipeline_dffe[13] (
	.clk(clock),
	.d(\op_1~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_13),
	.prn(vcc));
defparam \pipeline_dffe[13] .is_wysiwyg = "true";
defparam \pipeline_dffe[13] .power_up = "low";

dffeas \pipeline_dffe[12] (
	.clk(clock),
	.d(\op_1~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_12),
	.prn(vcc));
defparam \pipeline_dffe[12] .is_wysiwyg = "true";
defparam \pipeline_dffe[12] .power_up = "low";

dffeas \pipeline_dffe[11] (
	.clk(clock),
	.d(\op_1~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \pipeline_dffe[11] .is_wysiwyg = "true";
defparam \pipeline_dffe[11] .power_up = "low";

dffeas \pipeline_dffe[0] (
	.clk(clock),
	.d(\op_1~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_0),
	.prn(vcc));
defparam \pipeline_dffe[0] .is_wysiwyg = "true";
defparam \pipeline_dffe[0] .power_up = "low";

dffeas \pipeline_dffe[1] (
	.clk(clock),
	.d(\op_1~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_1),
	.prn(vcc));
defparam \pipeline_dffe[1] .is_wysiwyg = "true";
defparam \pipeline_dffe[1] .power_up = "low";

dffeas \pipeline_dffe[2] (
	.clk(clock),
	.d(\op_1~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \pipeline_dffe[2] .is_wysiwyg = "true";
defparam \pipeline_dffe[2] .power_up = "low";

dffeas \pipeline_dffe[3] (
	.clk(clock),
	.d(\op_1~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \pipeline_dffe[3] .is_wysiwyg = "true";
defparam \pipeline_dffe[3] .power_up = "low";

dffeas \pipeline_dffe[4] (
	.clk(clock),
	.d(\op_1~49_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \pipeline_dffe[4] .is_wysiwyg = "true";
defparam \pipeline_dffe[4] .power_up = "low";

dffeas \pipeline_dffe[5] (
	.clk(clock),
	.d(\op_1~53_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \pipeline_dffe[5] .is_wysiwyg = "true";
defparam \pipeline_dffe[5] .power_up = "low";

dffeas \pipeline_dffe[6] (
	.clk(clock),
	.d(\op_1~57_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \pipeline_dffe[6] .is_wysiwyg = "true";
defparam \pipeline_dffe[6] .power_up = "low";

dffeas \pipeline_dffe[7] (
	.clk(clock),
	.d(\op_1~61_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \pipeline_dffe[7] .is_wysiwyg = "true";
defparam \pipeline_dffe[7] .power_up = "low";

dffeas \pipeline_dffe[8] (
	.clk(clock),
	.d(\op_1~65_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \pipeline_dffe[8] .is_wysiwyg = "true";
defparam \pipeline_dffe[8] .power_up = "low";

dffeas \pipeline_dffe[9] (
	.clk(clock),
	.d(\op_1~69_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \pipeline_dffe[9] .is_wysiwyg = "true";
defparam \pipeline_dffe[9] .power_up = "low";

dffeas \pipeline_dffe[10] (
	.clk(clock),
	.d(\op_1~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \pipeline_dffe[10] .is_wysiwyg = "true";
defparam \pipeline_dffe[10] .power_up = "low";

arriav_lcell_comb \op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~29_sumout ),
	.cout(\op_1~30 ),
	.shareout());
defparam \op_1~29 .extended_lut = "off";
defparam \op_1~29 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~29 .shared_arith = "off";

arriav_lcell_comb \op_1~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_1),
	.datag(gnd),
	.cin(\op_1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~37_sumout ),
	.cout(\op_1~38 ),
	.shareout());
defparam \op_1~37 .extended_lut = "off";
defparam \op_1~37 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~37 .shared_arith = "off";

arriav_lcell_comb \op_1~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_2),
	.datag(gnd),
	.cin(\op_1~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~41_sumout ),
	.cout(\op_1~42 ),
	.shareout());
defparam \op_1~41 .extended_lut = "off";
defparam \op_1~41 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~41 .shared_arith = "off";

arriav_lcell_comb \op_1~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_3),
	.datag(gnd),
	.cin(\op_1~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~45_sumout ),
	.cout(\op_1~46 ),
	.shareout());
defparam \op_1~45 .extended_lut = "off";
defparam \op_1~45 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~45 .shared_arith = "off";

arriav_lcell_comb \op_1~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_4),
	.datag(gnd),
	.cin(\op_1~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~49_sumout ),
	.cout(\op_1~50 ),
	.shareout());
defparam \op_1~49 .extended_lut = "off";
defparam \op_1~49 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~49 .shared_arith = "off";

arriav_lcell_comb \op_1~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_5),
	.datag(gnd),
	.cin(\op_1~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~53_sumout ),
	.cout(\op_1~54 ),
	.shareout());
defparam \op_1~53 .extended_lut = "off";
defparam \op_1~53 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~53 .shared_arith = "off";

arriav_lcell_comb \op_1~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_6),
	.datag(gnd),
	.cin(\op_1~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~57_sumout ),
	.cout(\op_1~58 ),
	.shareout());
defparam \op_1~57 .extended_lut = "off";
defparam \op_1~57 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~57 .shared_arith = "off";

arriav_lcell_comb \op_1~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~61_sumout ),
	.cout(\op_1~62 ),
	.shareout());
defparam \op_1~61 .extended_lut = "off";
defparam \op_1~61 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~61 .shared_arith = "off";

arriav_lcell_comb \op_1~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~65_sumout ),
	.cout(\op_1~66 ),
	.shareout());
defparam \op_1~65 .extended_lut = "off";
defparam \op_1~65 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~65 .shared_arith = "off";

arriav_lcell_comb \op_1~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~69_sumout ),
	.cout(\op_1~70 ),
	.shareout());
defparam \op_1~69 .extended_lut = "off";
defparam \op_1~69 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~69 .shared_arith = "off";

arriav_lcell_comb \op_1~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~33_sumout ),
	.cout(\op_1~34 ),
	.shareout());
defparam \op_1~33 .extended_lut = "off";
defparam \op_1~33 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~33 .shared_arith = "off";

arriav_lcell_comb \op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~25_sumout ),
	.cout(\op_1~26 ),
	.shareout());
defparam \op_1~25 .extended_lut = "off";
defparam \op_1~25 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~25 .shared_arith = "off";

arriav_lcell_comb \op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~21_sumout ),
	.cout(\op_1~22 ),
	.shareout());
defparam \op_1~21 .extended_lut = "off";
defparam \op_1~21 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~21 .shared_arith = "off";

arriav_lcell_comb \op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~17_sumout ),
	.cout(\op_1~18 ),
	.shareout());
defparam \op_1~17 .extended_lut = "off";
defparam \op_1~17 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~17 .shared_arith = "off";

arriav_lcell_comb \op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~13_sumout ),
	.cout(\op_1~14 ),
	.shareout());
defparam \op_1~13 .extended_lut = "off";
defparam \op_1~13 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~13 .shared_arith = "off";

arriav_lcell_comb \op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~9_sumout ),
	.cout(\op_1~10 ),
	.shareout());
defparam \op_1~9 .extended_lut = "off";
defparam \op_1~9 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~9 .shared_arith = "off";

arriav_lcell_comb \op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_16),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~5_sumout ),
	.cout(\op_1~6 ),
	.shareout());
defparam \op_1~5 .extended_lut = "off";
defparam \op_1~5 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~5 .shared_arith = "off";

arriav_lcell_comb \op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_17),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~1_sumout ),
	.cout(),
	.shareout());
defparam \op_1~1 .extended_lut = "off";
defparam \op_1~1 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~1 .shared_arith = "off";

endmodule

module nco_test_cordic_axor_1p_lpm_8 (
	sin_o_0,
	pipeline_dffe_17,
	pipeline_dffe_16,
	dffe16,
	dffe18,
	pipeline_dffe_15,
	pipeline_dffe_171,
	pipeline_dffe_14,
	pipeline_dffe_161,
	pipeline_dffe_12,
	pipeline_dffe_13,
	dffe17,
	pipeline_dffe_0,
	pipeline_dffe_151,
	dffe161,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_141,
	dffe15,
	pipeline_dffe_131,
	dffe14,
	dffe12,
	dffe13,
	pipeline_dffe_121,
	pipeline_dffe_111,
	pipeline_dffe_01,
	pipeline_dffe_18,
	pipeline_dffe_21,
	pipeline_dffe_31,
	pipeline_dffe_41,
	pipeline_dffe_51,
	pipeline_dffe_61,
	pipeline_dffe_71,
	pipeline_dffe_81,
	pipeline_dffe_91,
	pipeline_dffe_101,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	sin_o_0;
output 	pipeline_dffe_17;
output 	pipeline_dffe_16;
input 	dffe16;
input 	dffe18;
output 	pipeline_dffe_15;
input 	pipeline_dffe_171;
output 	pipeline_dffe_14;
input 	pipeline_dffe_161;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
input 	dffe17;
output 	pipeline_dffe_0;
input 	pipeline_dffe_151;
input 	dffe161;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
input 	pipeline_dffe_141;
input 	dffe15;
input 	pipeline_dffe_131;
input 	dffe14;
input 	dffe12;
input 	dffe13;
input 	pipeline_dffe_121;
input 	pipeline_dffe_111;
input 	pipeline_dffe_01;
input 	pipeline_dffe_18;
input 	pipeline_dffe_21;
input 	pipeline_dffe_31;
input 	pipeline_dffe_41;
input 	pipeline_dffe_51;
input 	pipeline_dffe_61;
input 	pipeline_dffe_71;
input 	pipeline_dffe_81;
input 	pipeline_dffe_91;
input 	pipeline_dffe_101;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[17]~q ;
wire \xordvalue[10]~q ;
wire \Add0~1_sumout ;
wire \a[16]~q ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \a[15]~q ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \a[14]~q ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \a[13]~q ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \a[12]~q ;
wire \a[0]~q ;
wire \xordvalue[0]~q ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \a[11]~q ;
wire \a[1]~q ;
wire \xordvalue[1]~q ;
wire \a[2]~q ;
wire \xordvalue[2]~q ;
wire \a[3]~q ;
wire \xordvalue[3]~q ;
wire \a[4]~q ;
wire \xordvalue[4]~q ;
wire \a[5]~q ;
wire \xordvalue[5]~q ;
wire \a[6]~q ;
wire \a[7]~q ;
wire \a[8]~q ;
wire \a[9]~q ;
wire \a[10]~q ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~65_sumout ;
wire \Add0~66 ;
wire \Add0~69_sumout ;
wire \Add0~70 ;
wire \xordvalue~0_combout ;
wire \xordvalue~1_combout ;
wire \xordvalue~2_combout ;
wire \xordvalue~3_combout ;
wire \xordvalue~4_combout ;
wire \xordvalue~5_combout ;
wire \xordvalue~6_combout ;


nco_test_lpm_add_sub_10 u0(
	.a_17(\a[17]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.a_16(\a[16]~q ),
	.a_15(\a[15]~q ),
	.a_14(\a[14]~q ),
	.a_13(\a[13]~q ),
	.a_12(\a[12]~q ),
	.a_0(\a[0]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_11(\a[11]~q ),
	.a_1(\a[1]~q ),
	.xordvalue_1(\xordvalue[1]~q ),
	.a_2(\a[2]~q ),
	.xordvalue_2(\xordvalue[2]~q ),
	.a_3(\a[3]~q ),
	.xordvalue_3(\xordvalue[3]~q ),
	.a_4(\a[4]~q ),
	.xordvalue_4(\xordvalue[4]~q ),
	.a_5(\a[5]~q ),
	.xordvalue_5(\xordvalue[5]~q ),
	.a_6(\a[6]~q ),
	.a_7(\a[7]~q ),
	.a_8(\a[8]~q ),
	.a_9(\a[9]~q ),
	.a_10(\a[10]~q ),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[17] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[17]~q ),
	.prn(vcc));
defparam \a[17] .is_wysiwyg = "true";
defparam \a[17] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_171),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h00000000000000FF;
defparam \Add0~1 .shared_arith = "off";

dffeas \a[16] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[16]~q ),
	.prn(vcc));
defparam \a[16] .is_wysiwyg = "true";
defparam \a[16] .power_up = "low";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h00000000000000FF;
defparam \Add0~5 .shared_arith = "off";

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h00000000000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h00000000000000FF;
defparam \Add0~13 .shared_arith = "off";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h00000000000000FF;
defparam \Add0~17 .shared_arith = "off";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h00000000000000FF;
defparam \Add0~21 .shared_arith = "off";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \xordvalue[1] (
	.clk(clk),
	.d(\xordvalue~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[1]~q ),
	.prn(vcc));
defparam \xordvalue[1] .is_wysiwyg = "true";
defparam \xordvalue[1] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \xordvalue[2] (
	.clk(clk),
	.d(\xordvalue~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[2]~q ),
	.prn(vcc));
defparam \xordvalue[2] .is_wysiwyg = "true";
defparam \xordvalue[2] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \xordvalue[3] (
	.clk(clk),
	.d(\xordvalue~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[3]~q ),
	.prn(vcc));
defparam \xordvalue[3] .is_wysiwyg = "true";
defparam \xordvalue[3] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \xordvalue[4] (
	.clk(clk),
	.d(\xordvalue~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[4]~q ),
	.prn(vcc));
defparam \xordvalue[4] .is_wysiwyg = "true";
defparam \xordvalue[4] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \xordvalue[5] (
	.clk(clk),
	.d(\xordvalue~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[5]~q ),
	.prn(vcc));
defparam \xordvalue[5] .is_wysiwyg = "true";
defparam \xordvalue[5] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe16),
	.datae(gnd),
	.dataf(!pipeline_dffe_01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~25 .shared_arith = "off";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h00000000000000FF;
defparam \Add0~29 .shared_arith = "off";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_18),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h00000000000000FF;
defparam \Add0~33 .shared_arith = "off";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h00000000000000FF;
defparam \Add0~37 .shared_arith = "off";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h00000000000000FF;
defparam \Add0~41 .shared_arith = "off";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h00000000000000FF;
defparam \Add0~45 .shared_arith = "off";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout());
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h00000000000000FF;
defparam \Add0~49 .shared_arith = "off";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout());
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h00000000000000FF;
defparam \Add0~53 .shared_arith = "off";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout());
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h00000000000000FF;
defparam \Add0~57 .shared_arith = "off";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout());
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h00000000000000FF;
defparam \Add0~61 .shared_arith = "off";

arriav_lcell_comb \Add0~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~65_sumout ),
	.cout(\Add0~66 ),
	.shareout());
defparam \Add0~65 .extended_lut = "off";
defparam \Add0~65 .lut_mask = 64'h00000000000000FF;
defparam \Add0~65 .shared_arith = "off";

arriav_lcell_comb \Add0~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~69_sumout ),
	.cout(\Add0~70 ),
	.shareout());
defparam \Add0~69 .extended_lut = "off";
defparam \Add0~69 .lut_mask = 64'h00000000000000FF;
defparam \Add0~69 .shared_arith = "off";

arriav_lcell_comb \xordvalue~0 (
	.dataa(!dffe16),
	.datab(!dffe18),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

arriav_lcell_comb \xordvalue~1 (
	.dataa(!dffe16),
	.datab(!dffe12),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~1 .extended_lut = "off";
defparam \xordvalue~1 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~1 .shared_arith = "off";

arriav_lcell_comb \xordvalue~2 (
	.dataa(!dffe16),
	.datab(!dffe13),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~2 .extended_lut = "off";
defparam \xordvalue~2 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~2 .shared_arith = "off";

arriav_lcell_comb \xordvalue~3 (
	.dataa(!dffe16),
	.datab(!dffe14),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~3 .extended_lut = "off";
defparam \xordvalue~3 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~3 .shared_arith = "off";

arriav_lcell_comb \xordvalue~4 (
	.dataa(!dffe16),
	.datab(!dffe15),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~4 .extended_lut = "off";
defparam \xordvalue~4 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~4 .shared_arith = "off";

arriav_lcell_comb \xordvalue~5 (
	.dataa(!dffe16),
	.datab(!dffe161),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~5 .extended_lut = "off";
defparam \xordvalue~5 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~5 .shared_arith = "off";

arriav_lcell_comb \xordvalue~6 (
	.dataa(!dffe16),
	.datab(!dffe17),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~6 .extended_lut = "off";
defparam \xordvalue~6 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~6 .shared_arith = "off";

endmodule

module nco_test_lpm_add_sub_10 (
	a_17,
	xordvalue_10,
	a_16,
	a_15,
	a_14,
	a_13,
	a_12,
	a_0,
	xordvalue_0,
	a_11,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	a_4,
	xordvalue_4,
	a_5,
	xordvalue_5,
	a_6,
	a_7,
	a_8,
	a_9,
	a_10,
	pipeline_dffe_17,
	pipeline_dffe_16,
	pipeline_dffe_15,
	pipeline_dffe_14,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_10;
input 	a_16;
input 	a_15;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_0;
input 	xordvalue_0;
input 	a_11;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
input 	a_4;
input 	xordvalue_4;
input 	a_5;
input 	xordvalue_5;
input 	a_6;
input 	a_7;
input 	a_8;
input 	a_9;
input 	a_10;
output 	pipeline_dffe_17;
output 	pipeline_dffe_16;
output 	pipeline_dffe_15;
output 	pipeline_dffe_14;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_add_sub_0qg_8 auto_generated(
	.a_17(a_17),
	.xordvalue_10(xordvalue_10),
	.a_16(a_16),
	.a_15(a_15),
	.a_14(a_14),
	.a_13(a_13),
	.a_12(a_12),
	.a_0(a_0),
	.xordvalue_0(xordvalue_0),
	.a_11(a_11),
	.a_1(a_1),
	.xordvalue_1(xordvalue_1),
	.a_2(a_2),
	.xordvalue_2(xordvalue_2),
	.a_3(a_3),
	.xordvalue_3(xordvalue_3),
	.a_4(a_4),
	.xordvalue_4(xordvalue_4),
	.a_5(a_5),
	.xordvalue_5(xordvalue_5),
	.a_6(a_6),
	.a_7(a_7),
	.a_8(a_8),
	.a_9(a_9),
	.a_10(a_10),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module nco_test_add_sub_0qg_8 (
	a_17,
	xordvalue_10,
	a_16,
	a_15,
	a_14,
	a_13,
	a_12,
	a_0,
	xordvalue_0,
	a_11,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	a_4,
	xordvalue_4,
	a_5,
	xordvalue_5,
	a_6,
	a_7,
	a_8,
	a_9,
	a_10,
	pipeline_dffe_17,
	pipeline_dffe_16,
	pipeline_dffe_15,
	pipeline_dffe_14,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_10;
input 	a_16;
input 	a_15;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_0;
input 	xordvalue_0;
input 	a_11;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
input 	a_4;
input 	xordvalue_4;
input 	a_5;
input 	xordvalue_5;
input 	a_6;
input 	a_7;
input 	a_8;
input 	a_9;
input 	a_10;
output 	pipeline_dffe_17;
output 	pipeline_dffe_16;
output 	pipeline_dffe_15;
output 	pipeline_dffe_14;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \op_1~26 ;
wire \op_1~34 ;
wire \op_1~38 ;
wire \op_1~42 ;
wire \op_1~46 ;
wire \op_1~50 ;
wire \op_1~54 ;
wire \op_1~58 ;
wire \op_1~62 ;
wire \op_1~66 ;
wire \op_1~70 ;
wire \op_1~30 ;
wire \op_1~22 ;
wire \op_1~18 ;
wire \op_1~14 ;
wire \op_1~10 ;
wire \op_1~6 ;
wire \op_1~1_sumout ;
wire \op_1~5_sumout ;
wire \op_1~9_sumout ;
wire \op_1~13_sumout ;
wire \op_1~21_sumout ;
wire \op_1~17_sumout ;
wire \op_1~25_sumout ;
wire \op_1~33_sumout ;
wire \op_1~37_sumout ;
wire \op_1~41_sumout ;
wire \op_1~45_sumout ;
wire \op_1~49_sumout ;
wire \op_1~53_sumout ;
wire \op_1~57_sumout ;
wire \op_1~61_sumout ;
wire \op_1~65_sumout ;
wire \op_1~69_sumout ;
wire \op_1~29_sumout ;


dffeas \pipeline_dffe[17] (
	.clk(clock),
	.d(\op_1~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_17),
	.prn(vcc));
defparam \pipeline_dffe[17] .is_wysiwyg = "true";
defparam \pipeline_dffe[17] .power_up = "low";

dffeas \pipeline_dffe[16] (
	.clk(clock),
	.d(\op_1~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_16),
	.prn(vcc));
defparam \pipeline_dffe[16] .is_wysiwyg = "true";
defparam \pipeline_dffe[16] .power_up = "low";

dffeas \pipeline_dffe[15] (
	.clk(clock),
	.d(\op_1~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_15),
	.prn(vcc));
defparam \pipeline_dffe[15] .is_wysiwyg = "true";
defparam \pipeline_dffe[15] .power_up = "low";

dffeas \pipeline_dffe[14] (
	.clk(clock),
	.d(\op_1~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_14),
	.prn(vcc));
defparam \pipeline_dffe[14] .is_wysiwyg = "true";
defparam \pipeline_dffe[14] .power_up = "low";

dffeas \pipeline_dffe[12] (
	.clk(clock),
	.d(\op_1~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_12),
	.prn(vcc));
defparam \pipeline_dffe[12] .is_wysiwyg = "true";
defparam \pipeline_dffe[12] .power_up = "low";

dffeas \pipeline_dffe[13] (
	.clk(clock),
	.d(\op_1~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_13),
	.prn(vcc));
defparam \pipeline_dffe[13] .is_wysiwyg = "true";
defparam \pipeline_dffe[13] .power_up = "low";

dffeas \pipeline_dffe[0] (
	.clk(clock),
	.d(\op_1~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_0),
	.prn(vcc));
defparam \pipeline_dffe[0] .is_wysiwyg = "true";
defparam \pipeline_dffe[0] .power_up = "low";

dffeas \pipeline_dffe[1] (
	.clk(clock),
	.d(\op_1~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_1),
	.prn(vcc));
defparam \pipeline_dffe[1] .is_wysiwyg = "true";
defparam \pipeline_dffe[1] .power_up = "low";

dffeas \pipeline_dffe[2] (
	.clk(clock),
	.d(\op_1~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \pipeline_dffe[2] .is_wysiwyg = "true";
defparam \pipeline_dffe[2] .power_up = "low";

dffeas \pipeline_dffe[3] (
	.clk(clock),
	.d(\op_1~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \pipeline_dffe[3] .is_wysiwyg = "true";
defparam \pipeline_dffe[3] .power_up = "low";

dffeas \pipeline_dffe[4] (
	.clk(clock),
	.d(\op_1~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \pipeline_dffe[4] .is_wysiwyg = "true";
defparam \pipeline_dffe[4] .power_up = "low";

dffeas \pipeline_dffe[5] (
	.clk(clock),
	.d(\op_1~49_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \pipeline_dffe[5] .is_wysiwyg = "true";
defparam \pipeline_dffe[5] .power_up = "low";

dffeas \pipeline_dffe[6] (
	.clk(clock),
	.d(\op_1~53_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \pipeline_dffe[6] .is_wysiwyg = "true";
defparam \pipeline_dffe[6] .power_up = "low";

dffeas \pipeline_dffe[7] (
	.clk(clock),
	.d(\op_1~57_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \pipeline_dffe[7] .is_wysiwyg = "true";
defparam \pipeline_dffe[7] .power_up = "low";

dffeas \pipeline_dffe[8] (
	.clk(clock),
	.d(\op_1~61_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \pipeline_dffe[8] .is_wysiwyg = "true";
defparam \pipeline_dffe[8] .power_up = "low";

dffeas \pipeline_dffe[9] (
	.clk(clock),
	.d(\op_1~65_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \pipeline_dffe[9] .is_wysiwyg = "true";
defparam \pipeline_dffe[9] .power_up = "low";

dffeas \pipeline_dffe[10] (
	.clk(clock),
	.d(\op_1~69_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \pipeline_dffe[10] .is_wysiwyg = "true";
defparam \pipeline_dffe[10] .power_up = "low";

dffeas \pipeline_dffe[11] (
	.clk(clock),
	.d(\op_1~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \pipeline_dffe[11] .is_wysiwyg = "true";
defparam \pipeline_dffe[11] .power_up = "low";

arriav_lcell_comb \op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~25_sumout ),
	.cout(\op_1~26 ),
	.shareout());
defparam \op_1~25 .extended_lut = "off";
defparam \op_1~25 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~25 .shared_arith = "off";

arriav_lcell_comb \op_1~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_1),
	.datag(gnd),
	.cin(\op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~33_sumout ),
	.cout(\op_1~34 ),
	.shareout());
defparam \op_1~33 .extended_lut = "off";
defparam \op_1~33 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~33 .shared_arith = "off";

arriav_lcell_comb \op_1~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_2),
	.datag(gnd),
	.cin(\op_1~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~37_sumout ),
	.cout(\op_1~38 ),
	.shareout());
defparam \op_1~37 .extended_lut = "off";
defparam \op_1~37 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~37 .shared_arith = "off";

arriav_lcell_comb \op_1~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_3),
	.datag(gnd),
	.cin(\op_1~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~41_sumout ),
	.cout(\op_1~42 ),
	.shareout());
defparam \op_1~41 .extended_lut = "off";
defparam \op_1~41 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~41 .shared_arith = "off";

arriav_lcell_comb \op_1~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_4),
	.datag(gnd),
	.cin(\op_1~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~45_sumout ),
	.cout(\op_1~46 ),
	.shareout());
defparam \op_1~45 .extended_lut = "off";
defparam \op_1~45 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~45 .shared_arith = "off";

arriav_lcell_comb \op_1~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_5),
	.datag(gnd),
	.cin(\op_1~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~49_sumout ),
	.cout(\op_1~50 ),
	.shareout());
defparam \op_1~49 .extended_lut = "off";
defparam \op_1~49 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~49 .shared_arith = "off";

arriav_lcell_comb \op_1~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~53_sumout ),
	.cout(\op_1~54 ),
	.shareout());
defparam \op_1~53 .extended_lut = "off";
defparam \op_1~53 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~53 .shared_arith = "off";

arriav_lcell_comb \op_1~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~57_sumout ),
	.cout(\op_1~58 ),
	.shareout());
defparam \op_1~57 .extended_lut = "off";
defparam \op_1~57 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~57 .shared_arith = "off";

arriav_lcell_comb \op_1~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~61_sumout ),
	.cout(\op_1~62 ),
	.shareout());
defparam \op_1~61 .extended_lut = "off";
defparam \op_1~61 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~61 .shared_arith = "off";

arriav_lcell_comb \op_1~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~65_sumout ),
	.cout(\op_1~66 ),
	.shareout());
defparam \op_1~65 .extended_lut = "off";
defparam \op_1~65 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~65 .shared_arith = "off";

arriav_lcell_comb \op_1~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~69_sumout ),
	.cout(\op_1~70 ),
	.shareout());
defparam \op_1~69 .extended_lut = "off";
defparam \op_1~69 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~69 .shared_arith = "off";

arriav_lcell_comb \op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~29_sumout ),
	.cout(\op_1~30 ),
	.shareout());
defparam \op_1~29 .extended_lut = "off";
defparam \op_1~29 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~29 .shared_arith = "off";

arriav_lcell_comb \op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~21_sumout ),
	.cout(\op_1~22 ),
	.shareout());
defparam \op_1~21 .extended_lut = "off";
defparam \op_1~21 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~21 .shared_arith = "off";

arriav_lcell_comb \op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~17_sumout ),
	.cout(\op_1~18 ),
	.shareout());
defparam \op_1~17 .extended_lut = "off";
defparam \op_1~17 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~17 .shared_arith = "off";

arriav_lcell_comb \op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~13_sumout ),
	.cout(\op_1~14 ),
	.shareout());
defparam \op_1~13 .extended_lut = "off";
defparam \op_1~13 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~13 .shared_arith = "off";

arriav_lcell_comb \op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~9_sumout ),
	.cout(\op_1~10 ),
	.shareout());
defparam \op_1~9 .extended_lut = "off";
defparam \op_1~9 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~9 .shared_arith = "off";

arriav_lcell_comb \op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_16),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~5_sumout ),
	.cout(\op_1~6 ),
	.shareout());
defparam \op_1~5 .extended_lut = "off";
defparam \op_1~5 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~5 .shared_arith = "off";

arriav_lcell_comb \op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_17),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~1_sumout ),
	.cout(),
	.shareout());
defparam \op_1~1 .extended_lut = "off";
defparam \op_1~1 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~1 .shared_arith = "off";

endmodule

module nco_test_cordic_axor_1p_lpm_9 (
	sin_o_0,
	pipeline_dffe_17,
	pipeline_dffe_16,
	dffe16,
	pipeline_dffe_15,
	pipeline_dffe_171,
	dffe18,
	pipeline_dffe_14,
	pipeline_dffe_13,
	pipeline_dffe_0,
	dffe17,
	pipeline_dffe_161,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_12,
	dffe161,
	pipeline_dffe_151,
	dffe15,
	pipeline_dffe_141,
	dffe13,
	dffe14,
	pipeline_dffe_121,
	pipeline_dffe_131,
	pipeline_dffe_01,
	pipeline_dffe_18,
	pipeline_dffe_21,
	pipeline_dffe_31,
	pipeline_dffe_41,
	pipeline_dffe_51,
	pipeline_dffe_61,
	pipeline_dffe_71,
	pipeline_dffe_81,
	pipeline_dffe_91,
	pipeline_dffe_101,
	pipeline_dffe_111,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	sin_o_0;
output 	pipeline_dffe_17;
output 	pipeline_dffe_16;
input 	dffe16;
output 	pipeline_dffe_15;
input 	pipeline_dffe_171;
input 	dffe18;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
output 	pipeline_dffe_0;
input 	dffe17;
input 	pipeline_dffe_161;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
output 	pipeline_dffe_12;
input 	dffe161;
input 	pipeline_dffe_151;
input 	dffe15;
input 	pipeline_dffe_141;
input 	dffe13;
input 	dffe14;
input 	pipeline_dffe_121;
input 	pipeline_dffe_131;
input 	pipeline_dffe_01;
input 	pipeline_dffe_18;
input 	pipeline_dffe_21;
input 	pipeline_dffe_31;
input 	pipeline_dffe_41;
input 	pipeline_dffe_51;
input 	pipeline_dffe_61;
input 	pipeline_dffe_71;
input 	pipeline_dffe_81;
input 	pipeline_dffe_91;
input 	pipeline_dffe_101;
input 	pipeline_dffe_111;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[17]~q ;
wire \xordvalue[10]~q ;
wire \Add0~1_sumout ;
wire \a[16]~q ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \a[15]~q ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \a[14]~q ;
wire \a[13]~q ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \a[0]~q ;
wire \xordvalue[0]~q ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \a[12]~q ;
wire \a[1]~q ;
wire \xordvalue[1]~q ;
wire \a[2]~q ;
wire \xordvalue[2]~q ;
wire \a[3]~q ;
wire \xordvalue[3]~q ;
wire \a[4]~q ;
wire \xordvalue[4]~q ;
wire \a[5]~q ;
wire \a[6]~q ;
wire \a[7]~q ;
wire \a[8]~q ;
wire \a[9]~q ;
wire \a[10]~q ;
wire \a[11]~q ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~65_sumout ;
wire \Add0~66 ;
wire \Add0~69_sumout ;
wire \Add0~70 ;
wire \xordvalue~0_combout ;
wire \xordvalue~1_combout ;
wire \xordvalue~2_combout ;
wire \xordvalue~3_combout ;
wire \xordvalue~4_combout ;
wire \xordvalue~5_combout ;


nco_test_lpm_add_sub_11 u0(
	.a_17(\a[17]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.a_16(\a[16]~q ),
	.a_15(\a[15]~q ),
	.a_14(\a[14]~q ),
	.a_13(\a[13]~q ),
	.a_0(\a[0]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_12(\a[12]~q ),
	.a_1(\a[1]~q ),
	.xordvalue_1(\xordvalue[1]~q ),
	.a_2(\a[2]~q ),
	.xordvalue_2(\xordvalue[2]~q ),
	.a_3(\a[3]~q ),
	.xordvalue_3(\xordvalue[3]~q ),
	.a_4(\a[4]~q ),
	.xordvalue_4(\xordvalue[4]~q ),
	.a_5(\a[5]~q ),
	.a_6(\a[6]~q ),
	.a_7(\a[7]~q ),
	.a_8(\a[8]~q ),
	.a_9(\a[9]~q ),
	.a_10(\a[10]~q ),
	.a_11(\a[11]~q ),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_12(pipeline_dffe_12),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[17] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[17]~q ),
	.prn(vcc));
defparam \a[17] .is_wysiwyg = "true";
defparam \a[17] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_171),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h00000000000000FF;
defparam \Add0~1 .shared_arith = "off";

dffeas \a[16] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[16]~q ),
	.prn(vcc));
defparam \a[16] .is_wysiwyg = "true";
defparam \a[16] .power_up = "low";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h00000000000000FF;
defparam \Add0~5 .shared_arith = "off";

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h00000000000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h00000000000000FF;
defparam \Add0~13 .shared_arith = "off";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h00000000000000FF;
defparam \Add0~17 .shared_arith = "off";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \xordvalue[1] (
	.clk(clk),
	.d(\xordvalue~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[1]~q ),
	.prn(vcc));
defparam \xordvalue[1] .is_wysiwyg = "true";
defparam \xordvalue[1] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \xordvalue[2] (
	.clk(clk),
	.d(\xordvalue~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[2]~q ),
	.prn(vcc));
defparam \xordvalue[2] .is_wysiwyg = "true";
defparam \xordvalue[2] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \xordvalue[3] (
	.clk(clk),
	.d(\xordvalue~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[3]~q ),
	.prn(vcc));
defparam \xordvalue[3] .is_wysiwyg = "true";
defparam \xordvalue[3] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \xordvalue[4] (
	.clk(clk),
	.d(\xordvalue~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[4]~q ),
	.prn(vcc));
defparam \xordvalue[4] .is_wysiwyg = "true";
defparam \xordvalue[4] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe16),
	.datae(gnd),
	.dataf(!pipeline_dffe_01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~21 .shared_arith = "off";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h00000000000000FF;
defparam \Add0~25 .shared_arith = "off";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_18),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h00000000000000FF;
defparam \Add0~29 .shared_arith = "off";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h00000000000000FF;
defparam \Add0~33 .shared_arith = "off";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h00000000000000FF;
defparam \Add0~37 .shared_arith = "off";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h00000000000000FF;
defparam \Add0~41 .shared_arith = "off";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h00000000000000FF;
defparam \Add0~45 .shared_arith = "off";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout());
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h00000000000000FF;
defparam \Add0~49 .shared_arith = "off";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout());
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h00000000000000FF;
defparam \Add0~53 .shared_arith = "off";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout());
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h00000000000000FF;
defparam \Add0~57 .shared_arith = "off";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout());
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h00000000000000FF;
defparam \Add0~61 .shared_arith = "off";

arriav_lcell_comb \Add0~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~65_sumout ),
	.cout(\Add0~66 ),
	.shareout());
defparam \Add0~65 .extended_lut = "off";
defparam \Add0~65 .lut_mask = 64'h00000000000000FF;
defparam \Add0~65 .shared_arith = "off";

arriav_lcell_comb \Add0~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~69_sumout ),
	.cout(\Add0~70 ),
	.shareout());
defparam \Add0~69 .extended_lut = "off";
defparam \Add0~69 .lut_mask = 64'h00000000000000FF;
defparam \Add0~69 .shared_arith = "off";

arriav_lcell_comb \xordvalue~0 (
	.dataa(!dffe18),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

arriav_lcell_comb \xordvalue~1 (
	.dataa(!dffe13),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~1 .extended_lut = "off";
defparam \xordvalue~1 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~1 .shared_arith = "off";

arriav_lcell_comb \xordvalue~2 (
	.dataa(!dffe14),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~2 .extended_lut = "off";
defparam \xordvalue~2 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~2 .shared_arith = "off";

arriav_lcell_comb \xordvalue~3 (
	.dataa(!dffe15),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~3 .extended_lut = "off";
defparam \xordvalue~3 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~3 .shared_arith = "off";

arriav_lcell_comb \xordvalue~4 (
	.dataa(!dffe161),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~4 .extended_lut = "off";
defparam \xordvalue~4 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~4 .shared_arith = "off";

arriav_lcell_comb \xordvalue~5 (
	.dataa(!dffe17),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~5 .extended_lut = "off";
defparam \xordvalue~5 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~5 .shared_arith = "off";

endmodule

module nco_test_lpm_add_sub_11 (
	a_17,
	xordvalue_10,
	a_16,
	a_15,
	a_14,
	a_13,
	a_0,
	xordvalue_0,
	a_12,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	a_4,
	xordvalue_4,
	a_5,
	a_6,
	a_7,
	a_8,
	a_9,
	a_10,
	a_11,
	pipeline_dffe_17,
	pipeline_dffe_16,
	pipeline_dffe_15,
	pipeline_dffe_14,
	pipeline_dffe_13,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_12,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_10;
input 	a_16;
input 	a_15;
input 	a_14;
input 	a_13;
input 	a_0;
input 	xordvalue_0;
input 	a_12;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
input 	a_4;
input 	xordvalue_4;
input 	a_5;
input 	a_6;
input 	a_7;
input 	a_8;
input 	a_9;
input 	a_10;
input 	a_11;
output 	pipeline_dffe_17;
output 	pipeline_dffe_16;
output 	pipeline_dffe_15;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
output 	pipeline_dffe_12;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_add_sub_0qg_9 auto_generated(
	.a_17(a_17),
	.xordvalue_10(xordvalue_10),
	.a_16(a_16),
	.a_15(a_15),
	.a_14(a_14),
	.a_13(a_13),
	.a_0(a_0),
	.xordvalue_0(xordvalue_0),
	.a_12(a_12),
	.a_1(a_1),
	.xordvalue_1(xordvalue_1),
	.a_2(a_2),
	.xordvalue_2(xordvalue_2),
	.a_3(a_3),
	.xordvalue_3(xordvalue_3),
	.a_4(a_4),
	.xordvalue_4(xordvalue_4),
	.a_5(a_5),
	.a_6(a_6),
	.a_7(a_7),
	.a_8(a_8),
	.a_9(a_9),
	.a_10(a_10),
	.a_11(a_11),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_12(pipeline_dffe_12),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module nco_test_add_sub_0qg_9 (
	a_17,
	xordvalue_10,
	a_16,
	a_15,
	a_14,
	a_13,
	a_0,
	xordvalue_0,
	a_12,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	a_4,
	xordvalue_4,
	a_5,
	a_6,
	a_7,
	a_8,
	a_9,
	a_10,
	a_11,
	pipeline_dffe_17,
	pipeline_dffe_16,
	pipeline_dffe_15,
	pipeline_dffe_14,
	pipeline_dffe_13,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_12,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_10;
input 	a_16;
input 	a_15;
input 	a_14;
input 	a_13;
input 	a_0;
input 	xordvalue_0;
input 	a_12;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
input 	a_4;
input 	xordvalue_4;
input 	a_5;
input 	a_6;
input 	a_7;
input 	a_8;
input 	a_9;
input 	a_10;
input 	a_11;
output 	pipeline_dffe_17;
output 	pipeline_dffe_16;
output 	pipeline_dffe_15;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
output 	pipeline_dffe_12;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \op_1~22 ;
wire \op_1~30 ;
wire \op_1~34 ;
wire \op_1~38 ;
wire \op_1~42 ;
wire \op_1~46 ;
wire \op_1~50 ;
wire \op_1~54 ;
wire \op_1~58 ;
wire \op_1~62 ;
wire \op_1~66 ;
wire \op_1~70 ;
wire \op_1~26 ;
wire \op_1~18 ;
wire \op_1~14 ;
wire \op_1~10 ;
wire \op_1~6 ;
wire \op_1~1_sumout ;
wire \op_1~5_sumout ;
wire \op_1~9_sumout ;
wire \op_1~13_sumout ;
wire \op_1~17_sumout ;
wire \op_1~21_sumout ;
wire \op_1~29_sumout ;
wire \op_1~33_sumout ;
wire \op_1~37_sumout ;
wire \op_1~41_sumout ;
wire \op_1~45_sumout ;
wire \op_1~49_sumout ;
wire \op_1~53_sumout ;
wire \op_1~57_sumout ;
wire \op_1~61_sumout ;
wire \op_1~65_sumout ;
wire \op_1~69_sumout ;
wire \op_1~25_sumout ;


dffeas \pipeline_dffe[17] (
	.clk(clock),
	.d(\op_1~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_17),
	.prn(vcc));
defparam \pipeline_dffe[17] .is_wysiwyg = "true";
defparam \pipeline_dffe[17] .power_up = "low";

dffeas \pipeline_dffe[16] (
	.clk(clock),
	.d(\op_1~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_16),
	.prn(vcc));
defparam \pipeline_dffe[16] .is_wysiwyg = "true";
defparam \pipeline_dffe[16] .power_up = "low";

dffeas \pipeline_dffe[15] (
	.clk(clock),
	.d(\op_1~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_15),
	.prn(vcc));
defparam \pipeline_dffe[15] .is_wysiwyg = "true";
defparam \pipeline_dffe[15] .power_up = "low";

dffeas \pipeline_dffe[14] (
	.clk(clock),
	.d(\op_1~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_14),
	.prn(vcc));
defparam \pipeline_dffe[14] .is_wysiwyg = "true";
defparam \pipeline_dffe[14] .power_up = "low";

dffeas \pipeline_dffe[13] (
	.clk(clock),
	.d(\op_1~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_13),
	.prn(vcc));
defparam \pipeline_dffe[13] .is_wysiwyg = "true";
defparam \pipeline_dffe[13] .power_up = "low";

dffeas \pipeline_dffe[0] (
	.clk(clock),
	.d(\op_1~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_0),
	.prn(vcc));
defparam \pipeline_dffe[0] .is_wysiwyg = "true";
defparam \pipeline_dffe[0] .power_up = "low";

dffeas \pipeline_dffe[1] (
	.clk(clock),
	.d(\op_1~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_1),
	.prn(vcc));
defparam \pipeline_dffe[1] .is_wysiwyg = "true";
defparam \pipeline_dffe[1] .power_up = "low";

dffeas \pipeline_dffe[2] (
	.clk(clock),
	.d(\op_1~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \pipeline_dffe[2] .is_wysiwyg = "true";
defparam \pipeline_dffe[2] .power_up = "low";

dffeas \pipeline_dffe[3] (
	.clk(clock),
	.d(\op_1~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \pipeline_dffe[3] .is_wysiwyg = "true";
defparam \pipeline_dffe[3] .power_up = "low";

dffeas \pipeline_dffe[4] (
	.clk(clock),
	.d(\op_1~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \pipeline_dffe[4] .is_wysiwyg = "true";
defparam \pipeline_dffe[4] .power_up = "low";

dffeas \pipeline_dffe[5] (
	.clk(clock),
	.d(\op_1~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \pipeline_dffe[5] .is_wysiwyg = "true";
defparam \pipeline_dffe[5] .power_up = "low";

dffeas \pipeline_dffe[6] (
	.clk(clock),
	.d(\op_1~49_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \pipeline_dffe[6] .is_wysiwyg = "true";
defparam \pipeline_dffe[6] .power_up = "low";

dffeas \pipeline_dffe[7] (
	.clk(clock),
	.d(\op_1~53_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \pipeline_dffe[7] .is_wysiwyg = "true";
defparam \pipeline_dffe[7] .power_up = "low";

dffeas \pipeline_dffe[8] (
	.clk(clock),
	.d(\op_1~57_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \pipeline_dffe[8] .is_wysiwyg = "true";
defparam \pipeline_dffe[8] .power_up = "low";

dffeas \pipeline_dffe[9] (
	.clk(clock),
	.d(\op_1~61_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \pipeline_dffe[9] .is_wysiwyg = "true";
defparam \pipeline_dffe[9] .power_up = "low";

dffeas \pipeline_dffe[10] (
	.clk(clock),
	.d(\op_1~65_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \pipeline_dffe[10] .is_wysiwyg = "true";
defparam \pipeline_dffe[10] .power_up = "low";

dffeas \pipeline_dffe[11] (
	.clk(clock),
	.d(\op_1~69_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \pipeline_dffe[11] .is_wysiwyg = "true";
defparam \pipeline_dffe[11] .power_up = "low";

dffeas \pipeline_dffe[12] (
	.clk(clock),
	.d(\op_1~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_12),
	.prn(vcc));
defparam \pipeline_dffe[12] .is_wysiwyg = "true";
defparam \pipeline_dffe[12] .power_up = "low";

arriav_lcell_comb \op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~21_sumout ),
	.cout(\op_1~22 ),
	.shareout());
defparam \op_1~21 .extended_lut = "off";
defparam \op_1~21 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~21 .shared_arith = "off";

arriav_lcell_comb \op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_1),
	.datag(gnd),
	.cin(\op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~29_sumout ),
	.cout(\op_1~30 ),
	.shareout());
defparam \op_1~29 .extended_lut = "off";
defparam \op_1~29 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~29 .shared_arith = "off";

arriav_lcell_comb \op_1~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_2),
	.datag(gnd),
	.cin(\op_1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~33_sumout ),
	.cout(\op_1~34 ),
	.shareout());
defparam \op_1~33 .extended_lut = "off";
defparam \op_1~33 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~33 .shared_arith = "off";

arriav_lcell_comb \op_1~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_3),
	.datag(gnd),
	.cin(\op_1~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~37_sumout ),
	.cout(\op_1~38 ),
	.shareout());
defparam \op_1~37 .extended_lut = "off";
defparam \op_1~37 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~37 .shared_arith = "off";

arriav_lcell_comb \op_1~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_4),
	.datag(gnd),
	.cin(\op_1~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~41_sumout ),
	.cout(\op_1~42 ),
	.shareout());
defparam \op_1~41 .extended_lut = "off";
defparam \op_1~41 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~41 .shared_arith = "off";

arriav_lcell_comb \op_1~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~45_sumout ),
	.cout(\op_1~46 ),
	.shareout());
defparam \op_1~45 .extended_lut = "off";
defparam \op_1~45 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~45 .shared_arith = "off";

arriav_lcell_comb \op_1~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~49_sumout ),
	.cout(\op_1~50 ),
	.shareout());
defparam \op_1~49 .extended_lut = "off";
defparam \op_1~49 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~49 .shared_arith = "off";

arriav_lcell_comb \op_1~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~53_sumout ),
	.cout(\op_1~54 ),
	.shareout());
defparam \op_1~53 .extended_lut = "off";
defparam \op_1~53 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~53 .shared_arith = "off";

arriav_lcell_comb \op_1~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~57_sumout ),
	.cout(\op_1~58 ),
	.shareout());
defparam \op_1~57 .extended_lut = "off";
defparam \op_1~57 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~57 .shared_arith = "off";

arriav_lcell_comb \op_1~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~61_sumout ),
	.cout(\op_1~62 ),
	.shareout());
defparam \op_1~61 .extended_lut = "off";
defparam \op_1~61 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~61 .shared_arith = "off";

arriav_lcell_comb \op_1~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~65_sumout ),
	.cout(\op_1~66 ),
	.shareout());
defparam \op_1~65 .extended_lut = "off";
defparam \op_1~65 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~65 .shared_arith = "off";

arriav_lcell_comb \op_1~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~69_sumout ),
	.cout(\op_1~70 ),
	.shareout());
defparam \op_1~69 .extended_lut = "off";
defparam \op_1~69 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~69 .shared_arith = "off";

arriav_lcell_comb \op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~25_sumout ),
	.cout(\op_1~26 ),
	.shareout());
defparam \op_1~25 .extended_lut = "off";
defparam \op_1~25 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~25 .shared_arith = "off";

arriav_lcell_comb \op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~17_sumout ),
	.cout(\op_1~18 ),
	.shareout());
defparam \op_1~17 .extended_lut = "off";
defparam \op_1~17 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~17 .shared_arith = "off";

arriav_lcell_comb \op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~13_sumout ),
	.cout(\op_1~14 ),
	.shareout());
defparam \op_1~13 .extended_lut = "off";
defparam \op_1~13 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~13 .shared_arith = "off";

arriav_lcell_comb \op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~9_sumout ),
	.cout(\op_1~10 ),
	.shareout());
defparam \op_1~9 .extended_lut = "off";
defparam \op_1~9 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~9 .shared_arith = "off";

arriav_lcell_comb \op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_16),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~5_sumout ),
	.cout(\op_1~6 ),
	.shareout());
defparam \op_1~5 .extended_lut = "off";
defparam \op_1~5 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~5 .shared_arith = "off";

arriav_lcell_comb \op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_17),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~1_sumout ),
	.cout(),
	.shareout());
defparam \op_1~1 .extended_lut = "off";
defparam \op_1~1 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~1 .shared_arith = "off";

endmodule

module nco_test_cordic_axor_1p_lpm_10 (
	sin_o_0,
	pipeline_dffe_17,
	pipeline_dffe_16,
	dffe16,
	dffe18,
	pipeline_dffe_14,
	pipeline_dffe_15,
	pipeline_dffe_171,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_161,
	dffe17,
	pipeline_dffe_151,
	dffe161,
	dffe14,
	dffe15,
	pipeline_dffe_141,
	pipeline_dffe_131,
	pipeline_dffe_01,
	pipeline_dffe_18,
	pipeline_dffe_21,
	pipeline_dffe_31,
	pipeline_dffe_41,
	pipeline_dffe_51,
	pipeline_dffe_61,
	pipeline_dffe_71,
	pipeline_dffe_81,
	pipeline_dffe_91,
	pipeline_dffe_101,
	pipeline_dffe_111,
	pipeline_dffe_121,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	sin_o_0;
output 	pipeline_dffe_17;
output 	pipeline_dffe_16;
input 	dffe16;
input 	dffe18;
output 	pipeline_dffe_14;
output 	pipeline_dffe_15;
input 	pipeline_dffe_171;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
input 	pipeline_dffe_161;
input 	dffe17;
input 	pipeline_dffe_151;
input 	dffe161;
input 	dffe14;
input 	dffe15;
input 	pipeline_dffe_141;
input 	pipeline_dffe_131;
input 	pipeline_dffe_01;
input 	pipeline_dffe_18;
input 	pipeline_dffe_21;
input 	pipeline_dffe_31;
input 	pipeline_dffe_41;
input 	pipeline_dffe_51;
input 	pipeline_dffe_61;
input 	pipeline_dffe_71;
input 	pipeline_dffe_81;
input 	pipeline_dffe_91;
input 	pipeline_dffe_101;
input 	pipeline_dffe_111;
input 	pipeline_dffe_121;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[17]~q ;
wire \xordvalue[10]~q ;
wire \Add0~1_sumout ;
wire \a[16]~q ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \a[15]~q ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \a[14]~q ;
wire \a[0]~q ;
wire \xordvalue[0]~q ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \a[13]~q ;
wire \a[1]~q ;
wire \xordvalue[1]~q ;
wire \a[2]~q ;
wire \xordvalue[2]~q ;
wire \a[3]~q ;
wire \xordvalue[3]~q ;
wire \a[4]~q ;
wire \a[5]~q ;
wire \a[6]~q ;
wire \a[7]~q ;
wire \a[8]~q ;
wire \a[9]~q ;
wire \a[10]~q ;
wire \a[11]~q ;
wire \a[12]~q ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~65_sumout ;
wire \Add0~66 ;
wire \Add0~69_sumout ;
wire \Add0~70 ;
wire \xordvalue~0_combout ;
wire \xordvalue~1_combout ;
wire \xordvalue~2_combout ;
wire \xordvalue~3_combout ;
wire \xordvalue~4_combout ;


nco_test_lpm_add_sub_12 u0(
	.a_17(\a[17]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.a_16(\a[16]~q ),
	.a_15(\a[15]~q ),
	.a_14(\a[14]~q ),
	.a_0(\a[0]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_13(\a[13]~q ),
	.a_1(\a[1]~q ),
	.xordvalue_1(\xordvalue[1]~q ),
	.a_2(\a[2]~q ),
	.xordvalue_2(\xordvalue[2]~q ),
	.a_3(\a[3]~q ),
	.xordvalue_3(\xordvalue[3]~q ),
	.a_4(\a[4]~q ),
	.a_5(\a[5]~q ),
	.a_6(\a[6]~q ),
	.a_7(\a[7]~q ),
	.a_8(\a[8]~q ),
	.a_9(\a[9]~q ),
	.a_10(\a[10]~q ),
	.a_11(\a[11]~q ),
	.a_12(\a[12]~q ),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_13(pipeline_dffe_13),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[17] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[17]~q ),
	.prn(vcc));
defparam \a[17] .is_wysiwyg = "true";
defparam \a[17] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_171),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h00000000000000FF;
defparam \Add0~1 .shared_arith = "off";

dffeas \a[16] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[16]~q ),
	.prn(vcc));
defparam \a[16] .is_wysiwyg = "true";
defparam \a[16] .power_up = "low";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h00000000000000FF;
defparam \Add0~5 .shared_arith = "off";

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h00000000000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h00000000000000FF;
defparam \Add0~13 .shared_arith = "off";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \xordvalue[1] (
	.clk(clk),
	.d(\xordvalue~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[1]~q ),
	.prn(vcc));
defparam \xordvalue[1] .is_wysiwyg = "true";
defparam \xordvalue[1] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \xordvalue[2] (
	.clk(clk),
	.d(\xordvalue~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[2]~q ),
	.prn(vcc));
defparam \xordvalue[2] .is_wysiwyg = "true";
defparam \xordvalue[2] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \xordvalue[3] (
	.clk(clk),
	.d(\xordvalue~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[3]~q ),
	.prn(vcc));
defparam \xordvalue[3] .is_wysiwyg = "true";
defparam \xordvalue[3] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe16),
	.datae(gnd),
	.dataf(!pipeline_dffe_01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~17 .shared_arith = "off";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h00000000000000FF;
defparam \Add0~21 .shared_arith = "off";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_18),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h00000000000000FF;
defparam \Add0~25 .shared_arith = "off";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h00000000000000FF;
defparam \Add0~29 .shared_arith = "off";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h00000000000000FF;
defparam \Add0~33 .shared_arith = "off";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h00000000000000FF;
defparam \Add0~37 .shared_arith = "off";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h00000000000000FF;
defparam \Add0~41 .shared_arith = "off";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h00000000000000FF;
defparam \Add0~45 .shared_arith = "off";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout());
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h00000000000000FF;
defparam \Add0~49 .shared_arith = "off";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout());
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h00000000000000FF;
defparam \Add0~53 .shared_arith = "off";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout());
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h00000000000000FF;
defparam \Add0~57 .shared_arith = "off";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout());
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h00000000000000FF;
defparam \Add0~61 .shared_arith = "off";

arriav_lcell_comb \Add0~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~65_sumout ),
	.cout(\Add0~66 ),
	.shareout());
defparam \Add0~65 .extended_lut = "off";
defparam \Add0~65 .lut_mask = 64'h00000000000000FF;
defparam \Add0~65 .shared_arith = "off";

arriav_lcell_comb \Add0~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~69_sumout ),
	.cout(\Add0~70 ),
	.shareout());
defparam \Add0~69 .extended_lut = "off";
defparam \Add0~69 .lut_mask = 64'h00000000000000FF;
defparam \Add0~69 .shared_arith = "off";

arriav_lcell_comb \xordvalue~0 (
	.dataa(!dffe16),
	.datab(!dffe18),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

arriav_lcell_comb \xordvalue~1 (
	.dataa(!dffe16),
	.datab(!dffe14),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~1 .extended_lut = "off";
defparam \xordvalue~1 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~1 .shared_arith = "off";

arriav_lcell_comb \xordvalue~2 (
	.dataa(!dffe16),
	.datab(!dffe15),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~2 .extended_lut = "off";
defparam \xordvalue~2 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~2 .shared_arith = "off";

arriav_lcell_comb \xordvalue~3 (
	.dataa(!dffe16),
	.datab(!dffe161),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~3 .extended_lut = "off";
defparam \xordvalue~3 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~3 .shared_arith = "off";

arriav_lcell_comb \xordvalue~4 (
	.dataa(!dffe16),
	.datab(!dffe17),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~4 .extended_lut = "off";
defparam \xordvalue~4 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~4 .shared_arith = "off";

endmodule

module nco_test_lpm_add_sub_12 (
	a_17,
	xordvalue_10,
	a_16,
	a_15,
	a_14,
	a_0,
	xordvalue_0,
	a_13,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	a_4,
	a_5,
	a_6,
	a_7,
	a_8,
	a_9,
	a_10,
	a_11,
	a_12,
	pipeline_dffe_17,
	pipeline_dffe_16,
	pipeline_dffe_14,
	pipeline_dffe_15,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_12,
	pipeline_dffe_13,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_10;
input 	a_16;
input 	a_15;
input 	a_14;
input 	a_0;
input 	xordvalue_0;
input 	a_13;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
input 	a_4;
input 	a_5;
input 	a_6;
input 	a_7;
input 	a_8;
input 	a_9;
input 	a_10;
input 	a_11;
input 	a_12;
output 	pipeline_dffe_17;
output 	pipeline_dffe_16;
output 	pipeline_dffe_14;
output 	pipeline_dffe_15;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_add_sub_0qg_10 auto_generated(
	.a_17(a_17),
	.xordvalue_10(xordvalue_10),
	.a_16(a_16),
	.a_15(a_15),
	.a_14(a_14),
	.a_0(a_0),
	.xordvalue_0(xordvalue_0),
	.a_13(a_13),
	.a_1(a_1),
	.xordvalue_1(xordvalue_1),
	.a_2(a_2),
	.xordvalue_2(xordvalue_2),
	.a_3(a_3),
	.xordvalue_3(xordvalue_3),
	.a_4(a_4),
	.a_5(a_5),
	.a_6(a_6),
	.a_7(a_7),
	.a_8(a_8),
	.a_9(a_9),
	.a_10(a_10),
	.a_11(a_11),
	.a_12(a_12),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_13(pipeline_dffe_13),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module nco_test_add_sub_0qg_10 (
	a_17,
	xordvalue_10,
	a_16,
	a_15,
	a_14,
	a_0,
	xordvalue_0,
	a_13,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	a_4,
	a_5,
	a_6,
	a_7,
	a_8,
	a_9,
	a_10,
	a_11,
	a_12,
	pipeline_dffe_17,
	pipeline_dffe_16,
	pipeline_dffe_14,
	pipeline_dffe_15,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_12,
	pipeline_dffe_13,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_10;
input 	a_16;
input 	a_15;
input 	a_14;
input 	a_0;
input 	xordvalue_0;
input 	a_13;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
input 	a_4;
input 	a_5;
input 	a_6;
input 	a_7;
input 	a_8;
input 	a_9;
input 	a_10;
input 	a_11;
input 	a_12;
output 	pipeline_dffe_17;
output 	pipeline_dffe_16;
output 	pipeline_dffe_14;
output 	pipeline_dffe_15;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \op_1~18 ;
wire \op_1~26 ;
wire \op_1~30 ;
wire \op_1~34 ;
wire \op_1~38 ;
wire \op_1~42 ;
wire \op_1~46 ;
wire \op_1~50 ;
wire \op_1~54 ;
wire \op_1~58 ;
wire \op_1~62 ;
wire \op_1~66 ;
wire \op_1~70 ;
wire \op_1~22 ;
wire \op_1~14 ;
wire \op_1~10 ;
wire \op_1~6 ;
wire \op_1~1_sumout ;
wire \op_1~5_sumout ;
wire \op_1~13_sumout ;
wire \op_1~9_sumout ;
wire \op_1~17_sumout ;
wire \op_1~25_sumout ;
wire \op_1~29_sumout ;
wire \op_1~33_sumout ;
wire \op_1~37_sumout ;
wire \op_1~41_sumout ;
wire \op_1~45_sumout ;
wire \op_1~49_sumout ;
wire \op_1~53_sumout ;
wire \op_1~57_sumout ;
wire \op_1~61_sumout ;
wire \op_1~65_sumout ;
wire \op_1~69_sumout ;
wire \op_1~21_sumout ;


dffeas \pipeline_dffe[17] (
	.clk(clock),
	.d(\op_1~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_17),
	.prn(vcc));
defparam \pipeline_dffe[17] .is_wysiwyg = "true";
defparam \pipeline_dffe[17] .power_up = "low";

dffeas \pipeline_dffe[16] (
	.clk(clock),
	.d(\op_1~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_16),
	.prn(vcc));
defparam \pipeline_dffe[16] .is_wysiwyg = "true";
defparam \pipeline_dffe[16] .power_up = "low";

dffeas \pipeline_dffe[14] (
	.clk(clock),
	.d(\op_1~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_14),
	.prn(vcc));
defparam \pipeline_dffe[14] .is_wysiwyg = "true";
defparam \pipeline_dffe[14] .power_up = "low";

dffeas \pipeline_dffe[15] (
	.clk(clock),
	.d(\op_1~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_15),
	.prn(vcc));
defparam \pipeline_dffe[15] .is_wysiwyg = "true";
defparam \pipeline_dffe[15] .power_up = "low";

dffeas \pipeline_dffe[0] (
	.clk(clock),
	.d(\op_1~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_0),
	.prn(vcc));
defparam \pipeline_dffe[0] .is_wysiwyg = "true";
defparam \pipeline_dffe[0] .power_up = "low";

dffeas \pipeline_dffe[1] (
	.clk(clock),
	.d(\op_1~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_1),
	.prn(vcc));
defparam \pipeline_dffe[1] .is_wysiwyg = "true";
defparam \pipeline_dffe[1] .power_up = "low";

dffeas \pipeline_dffe[2] (
	.clk(clock),
	.d(\op_1~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \pipeline_dffe[2] .is_wysiwyg = "true";
defparam \pipeline_dffe[2] .power_up = "low";

dffeas \pipeline_dffe[3] (
	.clk(clock),
	.d(\op_1~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \pipeline_dffe[3] .is_wysiwyg = "true";
defparam \pipeline_dffe[3] .power_up = "low";

dffeas \pipeline_dffe[4] (
	.clk(clock),
	.d(\op_1~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \pipeline_dffe[4] .is_wysiwyg = "true";
defparam \pipeline_dffe[4] .power_up = "low";

dffeas \pipeline_dffe[5] (
	.clk(clock),
	.d(\op_1~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \pipeline_dffe[5] .is_wysiwyg = "true";
defparam \pipeline_dffe[5] .power_up = "low";

dffeas \pipeline_dffe[6] (
	.clk(clock),
	.d(\op_1~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \pipeline_dffe[6] .is_wysiwyg = "true";
defparam \pipeline_dffe[6] .power_up = "low";

dffeas \pipeline_dffe[7] (
	.clk(clock),
	.d(\op_1~49_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \pipeline_dffe[7] .is_wysiwyg = "true";
defparam \pipeline_dffe[7] .power_up = "low";

dffeas \pipeline_dffe[8] (
	.clk(clock),
	.d(\op_1~53_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \pipeline_dffe[8] .is_wysiwyg = "true";
defparam \pipeline_dffe[8] .power_up = "low";

dffeas \pipeline_dffe[9] (
	.clk(clock),
	.d(\op_1~57_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \pipeline_dffe[9] .is_wysiwyg = "true";
defparam \pipeline_dffe[9] .power_up = "low";

dffeas \pipeline_dffe[10] (
	.clk(clock),
	.d(\op_1~61_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \pipeline_dffe[10] .is_wysiwyg = "true";
defparam \pipeline_dffe[10] .power_up = "low";

dffeas \pipeline_dffe[11] (
	.clk(clock),
	.d(\op_1~65_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \pipeline_dffe[11] .is_wysiwyg = "true";
defparam \pipeline_dffe[11] .power_up = "low";

dffeas \pipeline_dffe[12] (
	.clk(clock),
	.d(\op_1~69_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_12),
	.prn(vcc));
defparam \pipeline_dffe[12] .is_wysiwyg = "true";
defparam \pipeline_dffe[12] .power_up = "low";

dffeas \pipeline_dffe[13] (
	.clk(clock),
	.d(\op_1~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_13),
	.prn(vcc));
defparam \pipeline_dffe[13] .is_wysiwyg = "true";
defparam \pipeline_dffe[13] .power_up = "low";

arriav_lcell_comb \op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~17_sumout ),
	.cout(\op_1~18 ),
	.shareout());
defparam \op_1~17 .extended_lut = "off";
defparam \op_1~17 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~17 .shared_arith = "off";

arriav_lcell_comb \op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_1),
	.datag(gnd),
	.cin(\op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~25_sumout ),
	.cout(\op_1~26 ),
	.shareout());
defparam \op_1~25 .extended_lut = "off";
defparam \op_1~25 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~25 .shared_arith = "off";

arriav_lcell_comb \op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_2),
	.datag(gnd),
	.cin(\op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~29_sumout ),
	.cout(\op_1~30 ),
	.shareout());
defparam \op_1~29 .extended_lut = "off";
defparam \op_1~29 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~29 .shared_arith = "off";

arriav_lcell_comb \op_1~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_3),
	.datag(gnd),
	.cin(\op_1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~33_sumout ),
	.cout(\op_1~34 ),
	.shareout());
defparam \op_1~33 .extended_lut = "off";
defparam \op_1~33 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~33 .shared_arith = "off";

arriav_lcell_comb \op_1~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~37_sumout ),
	.cout(\op_1~38 ),
	.shareout());
defparam \op_1~37 .extended_lut = "off";
defparam \op_1~37 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~37 .shared_arith = "off";

arriav_lcell_comb \op_1~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~41_sumout ),
	.cout(\op_1~42 ),
	.shareout());
defparam \op_1~41 .extended_lut = "off";
defparam \op_1~41 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~41 .shared_arith = "off";

arriav_lcell_comb \op_1~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~45_sumout ),
	.cout(\op_1~46 ),
	.shareout());
defparam \op_1~45 .extended_lut = "off";
defparam \op_1~45 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~45 .shared_arith = "off";

arriav_lcell_comb \op_1~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~49_sumout ),
	.cout(\op_1~50 ),
	.shareout());
defparam \op_1~49 .extended_lut = "off";
defparam \op_1~49 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~49 .shared_arith = "off";

arriav_lcell_comb \op_1~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~53_sumout ),
	.cout(\op_1~54 ),
	.shareout());
defparam \op_1~53 .extended_lut = "off";
defparam \op_1~53 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~53 .shared_arith = "off";

arriav_lcell_comb \op_1~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~57_sumout ),
	.cout(\op_1~58 ),
	.shareout());
defparam \op_1~57 .extended_lut = "off";
defparam \op_1~57 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~57 .shared_arith = "off";

arriav_lcell_comb \op_1~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~61_sumout ),
	.cout(\op_1~62 ),
	.shareout());
defparam \op_1~61 .extended_lut = "off";
defparam \op_1~61 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~61 .shared_arith = "off";

arriav_lcell_comb \op_1~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~65_sumout ),
	.cout(\op_1~66 ),
	.shareout());
defparam \op_1~65 .extended_lut = "off";
defparam \op_1~65 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~65 .shared_arith = "off";

arriav_lcell_comb \op_1~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~69_sumout ),
	.cout(\op_1~70 ),
	.shareout());
defparam \op_1~69 .extended_lut = "off";
defparam \op_1~69 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~69 .shared_arith = "off";

arriav_lcell_comb \op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~21_sumout ),
	.cout(\op_1~22 ),
	.shareout());
defparam \op_1~21 .extended_lut = "off";
defparam \op_1~21 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~21 .shared_arith = "off";

arriav_lcell_comb \op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~13_sumout ),
	.cout(\op_1~14 ),
	.shareout());
defparam \op_1~13 .extended_lut = "off";
defparam \op_1~13 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~13 .shared_arith = "off";

arriav_lcell_comb \op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~9_sumout ),
	.cout(\op_1~10 ),
	.shareout());
defparam \op_1~9 .extended_lut = "off";
defparam \op_1~9 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~9 .shared_arith = "off";

arriav_lcell_comb \op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_16),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~5_sumout ),
	.cout(\op_1~6 ),
	.shareout());
defparam \op_1~5 .extended_lut = "off";
defparam \op_1~5 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~5 .shared_arith = "off";

arriav_lcell_comb \op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_17),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~1_sumout ),
	.cout(),
	.shareout());
defparam \op_1~1 .extended_lut = "off";
defparam \op_1~1 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~1 .shared_arith = "off";

endmodule

module nco_test_cordic_axor_1p_lpm_11 (
	sin_o_0,
	pipeline_dffe_17,
	pipeline_dffe_16,
	pipeline_dffe_15,
	pipeline_dffe_0,
	dffe16,
	pipeline_dffe_171,
	dffe18,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	dffe17,
	pipeline_dffe_161,
	dffe15,
	dffe161,
	pipeline_dffe_141,
	pipeline_dffe_151,
	pipeline_dffe_01,
	pipeline_dffe_18,
	pipeline_dffe_21,
	pipeline_dffe_31,
	pipeline_dffe_41,
	pipeline_dffe_51,
	pipeline_dffe_61,
	pipeline_dffe_71,
	pipeline_dffe_81,
	pipeline_dffe_91,
	pipeline_dffe_101,
	pipeline_dffe_111,
	pipeline_dffe_121,
	pipeline_dffe_131,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	sin_o_0;
output 	pipeline_dffe_17;
output 	pipeline_dffe_16;
output 	pipeline_dffe_15;
output 	pipeline_dffe_0;
input 	dffe16;
input 	pipeline_dffe_171;
input 	dffe18;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
input 	dffe17;
input 	pipeline_dffe_161;
input 	dffe15;
input 	dffe161;
input 	pipeline_dffe_141;
input 	pipeline_dffe_151;
input 	pipeline_dffe_01;
input 	pipeline_dffe_18;
input 	pipeline_dffe_21;
input 	pipeline_dffe_31;
input 	pipeline_dffe_41;
input 	pipeline_dffe_51;
input 	pipeline_dffe_61;
input 	pipeline_dffe_71;
input 	pipeline_dffe_81;
input 	pipeline_dffe_91;
input 	pipeline_dffe_101;
input 	pipeline_dffe_111;
input 	pipeline_dffe_121;
input 	pipeline_dffe_131;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[17]~q ;
wire \xordvalue[10]~q ;
wire \Add0~1_sumout ;
wire \a[16]~q ;
wire \a[15]~q ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \a[0]~q ;
wire \xordvalue[0]~q ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \a[14]~q ;
wire \a[1]~q ;
wire \xordvalue[1]~q ;
wire \a[2]~q ;
wire \xordvalue[2]~q ;
wire \a[3]~q ;
wire \a[4]~q ;
wire \a[5]~q ;
wire \a[6]~q ;
wire \a[7]~q ;
wire \a[8]~q ;
wire \a[9]~q ;
wire \a[10]~q ;
wire \a[11]~q ;
wire \a[12]~q ;
wire \a[13]~q ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~65_sumout ;
wire \Add0~66 ;
wire \Add0~69_sumout ;
wire \Add0~70 ;
wire \xordvalue~0_combout ;
wire \xordvalue~1_combout ;
wire \xordvalue~2_combout ;
wire \xordvalue~3_combout ;


nco_test_lpm_add_sub_13 u0(
	.a_17(\a[17]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.a_16(\a[16]~q ),
	.a_15(\a[15]~q ),
	.a_0(\a[0]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_14(\a[14]~q ),
	.a_1(\a[1]~q ),
	.xordvalue_1(\xordvalue[1]~q ),
	.a_2(\a[2]~q ),
	.xordvalue_2(\xordvalue[2]~q ),
	.a_3(\a[3]~q ),
	.a_4(\a[4]~q ),
	.a_5(\a[5]~q ),
	.a_6(\a[6]~q ),
	.a_7(\a[7]~q ),
	.a_8(\a[8]~q ),
	.a_9(\a[9]~q ),
	.a_10(\a[10]~q ),
	.a_11(\a[11]~q ),
	.a_12(\a[12]~q ),
	.a_13(\a[13]~q ),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_14(pipeline_dffe_14),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[17] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[17]~q ),
	.prn(vcc));
defparam \a[17] .is_wysiwyg = "true";
defparam \a[17] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_171),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h00000000000000FF;
defparam \Add0~1 .shared_arith = "off";

dffeas \a[16] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[16]~q ),
	.prn(vcc));
defparam \a[16] .is_wysiwyg = "true";
defparam \a[16] .power_up = "low";

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h00000000000000FF;
defparam \Add0~5 .shared_arith = "off";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h00000000000000FF;
defparam \Add0~9 .shared_arith = "off";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \xordvalue[1] (
	.clk(clk),
	.d(\xordvalue~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[1]~q ),
	.prn(vcc));
defparam \xordvalue[1] .is_wysiwyg = "true";
defparam \xordvalue[1] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \xordvalue[2] (
	.clk(clk),
	.d(\xordvalue~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[2]~q ),
	.prn(vcc));
defparam \xordvalue[2] .is_wysiwyg = "true";
defparam \xordvalue[2] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe16),
	.datae(gnd),
	.dataf(!pipeline_dffe_01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~13 .shared_arith = "off";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h00000000000000FF;
defparam \Add0~17 .shared_arith = "off";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_18),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h00000000000000FF;
defparam \Add0~21 .shared_arith = "off";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h00000000000000FF;
defparam \Add0~25 .shared_arith = "off";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h00000000000000FF;
defparam \Add0~29 .shared_arith = "off";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h00000000000000FF;
defparam \Add0~33 .shared_arith = "off";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h00000000000000FF;
defparam \Add0~37 .shared_arith = "off";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h00000000000000FF;
defparam \Add0~41 .shared_arith = "off";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h00000000000000FF;
defparam \Add0~45 .shared_arith = "off";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout());
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h00000000000000FF;
defparam \Add0~49 .shared_arith = "off";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout());
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h00000000000000FF;
defparam \Add0~53 .shared_arith = "off";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout());
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h00000000000000FF;
defparam \Add0~57 .shared_arith = "off";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout());
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h00000000000000FF;
defparam \Add0~61 .shared_arith = "off";

arriav_lcell_comb \Add0~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~65_sumout ),
	.cout(\Add0~66 ),
	.shareout());
defparam \Add0~65 .extended_lut = "off";
defparam \Add0~65 .lut_mask = 64'h00000000000000FF;
defparam \Add0~65 .shared_arith = "off";

arriav_lcell_comb \Add0~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~69_sumout ),
	.cout(\Add0~70 ),
	.shareout());
defparam \Add0~69 .extended_lut = "off";
defparam \Add0~69 .lut_mask = 64'h00000000000000FF;
defparam \Add0~69 .shared_arith = "off";

arriav_lcell_comb \xordvalue~0 (
	.dataa(!dffe18),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

arriav_lcell_comb \xordvalue~1 (
	.dataa(!dffe15),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~1 .extended_lut = "off";
defparam \xordvalue~1 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~1 .shared_arith = "off";

arriav_lcell_comb \xordvalue~2 (
	.dataa(!dffe161),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~2 .extended_lut = "off";
defparam \xordvalue~2 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~2 .shared_arith = "off";

arriav_lcell_comb \xordvalue~3 (
	.dataa(!dffe17),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~3 .extended_lut = "off";
defparam \xordvalue~3 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~3 .shared_arith = "off";

endmodule

module nco_test_lpm_add_sub_13 (
	a_17,
	xordvalue_10,
	a_16,
	a_15,
	a_0,
	xordvalue_0,
	a_14,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	a_4,
	a_5,
	a_6,
	a_7,
	a_8,
	a_9,
	a_10,
	a_11,
	a_12,
	a_13,
	pipeline_dffe_17,
	pipeline_dffe_16,
	pipeline_dffe_15,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_10;
input 	a_16;
input 	a_15;
input 	a_0;
input 	xordvalue_0;
input 	a_14;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	a_4;
input 	a_5;
input 	a_6;
input 	a_7;
input 	a_8;
input 	a_9;
input 	a_10;
input 	a_11;
input 	a_12;
input 	a_13;
output 	pipeline_dffe_17;
output 	pipeline_dffe_16;
output 	pipeline_dffe_15;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_add_sub_0qg_11 auto_generated(
	.a_17(a_17),
	.xordvalue_10(xordvalue_10),
	.a_16(a_16),
	.a_15(a_15),
	.a_0(a_0),
	.xordvalue_0(xordvalue_0),
	.a_14(a_14),
	.a_1(a_1),
	.xordvalue_1(xordvalue_1),
	.a_2(a_2),
	.xordvalue_2(xordvalue_2),
	.a_3(a_3),
	.a_4(a_4),
	.a_5(a_5),
	.a_6(a_6),
	.a_7(a_7),
	.a_8(a_8),
	.a_9(a_9),
	.a_10(a_10),
	.a_11(a_11),
	.a_12(a_12),
	.a_13(a_13),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_14(pipeline_dffe_14),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module nco_test_add_sub_0qg_11 (
	a_17,
	xordvalue_10,
	a_16,
	a_15,
	a_0,
	xordvalue_0,
	a_14,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	a_4,
	a_5,
	a_6,
	a_7,
	a_8,
	a_9,
	a_10,
	a_11,
	a_12,
	a_13,
	pipeline_dffe_17,
	pipeline_dffe_16,
	pipeline_dffe_15,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_10;
input 	a_16;
input 	a_15;
input 	a_0;
input 	xordvalue_0;
input 	a_14;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	a_4;
input 	a_5;
input 	a_6;
input 	a_7;
input 	a_8;
input 	a_9;
input 	a_10;
input 	a_11;
input 	a_12;
input 	a_13;
output 	pipeline_dffe_17;
output 	pipeline_dffe_16;
output 	pipeline_dffe_15;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \op_1~14 ;
wire \op_1~22 ;
wire \op_1~26 ;
wire \op_1~30 ;
wire \op_1~34 ;
wire \op_1~38 ;
wire \op_1~42 ;
wire \op_1~46 ;
wire \op_1~50 ;
wire \op_1~54 ;
wire \op_1~58 ;
wire \op_1~62 ;
wire \op_1~66 ;
wire \op_1~70 ;
wire \op_1~18 ;
wire \op_1~10 ;
wire \op_1~6 ;
wire \op_1~1_sumout ;
wire \op_1~5_sumout ;
wire \op_1~9_sumout ;
wire \op_1~13_sumout ;
wire \op_1~21_sumout ;
wire \op_1~25_sumout ;
wire \op_1~29_sumout ;
wire \op_1~33_sumout ;
wire \op_1~37_sumout ;
wire \op_1~41_sumout ;
wire \op_1~45_sumout ;
wire \op_1~49_sumout ;
wire \op_1~53_sumout ;
wire \op_1~57_sumout ;
wire \op_1~61_sumout ;
wire \op_1~65_sumout ;
wire \op_1~69_sumout ;
wire \op_1~17_sumout ;


dffeas \pipeline_dffe[17] (
	.clk(clock),
	.d(\op_1~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_17),
	.prn(vcc));
defparam \pipeline_dffe[17] .is_wysiwyg = "true";
defparam \pipeline_dffe[17] .power_up = "low";

dffeas \pipeline_dffe[16] (
	.clk(clock),
	.d(\op_1~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_16),
	.prn(vcc));
defparam \pipeline_dffe[16] .is_wysiwyg = "true";
defparam \pipeline_dffe[16] .power_up = "low";

dffeas \pipeline_dffe[15] (
	.clk(clock),
	.d(\op_1~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_15),
	.prn(vcc));
defparam \pipeline_dffe[15] .is_wysiwyg = "true";
defparam \pipeline_dffe[15] .power_up = "low";

dffeas \pipeline_dffe[0] (
	.clk(clock),
	.d(\op_1~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_0),
	.prn(vcc));
defparam \pipeline_dffe[0] .is_wysiwyg = "true";
defparam \pipeline_dffe[0] .power_up = "low";

dffeas \pipeline_dffe[1] (
	.clk(clock),
	.d(\op_1~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_1),
	.prn(vcc));
defparam \pipeline_dffe[1] .is_wysiwyg = "true";
defparam \pipeline_dffe[1] .power_up = "low";

dffeas \pipeline_dffe[2] (
	.clk(clock),
	.d(\op_1~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \pipeline_dffe[2] .is_wysiwyg = "true";
defparam \pipeline_dffe[2] .power_up = "low";

dffeas \pipeline_dffe[3] (
	.clk(clock),
	.d(\op_1~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \pipeline_dffe[3] .is_wysiwyg = "true";
defparam \pipeline_dffe[3] .power_up = "low";

dffeas \pipeline_dffe[4] (
	.clk(clock),
	.d(\op_1~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \pipeline_dffe[4] .is_wysiwyg = "true";
defparam \pipeline_dffe[4] .power_up = "low";

dffeas \pipeline_dffe[5] (
	.clk(clock),
	.d(\op_1~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \pipeline_dffe[5] .is_wysiwyg = "true";
defparam \pipeline_dffe[5] .power_up = "low";

dffeas \pipeline_dffe[6] (
	.clk(clock),
	.d(\op_1~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \pipeline_dffe[6] .is_wysiwyg = "true";
defparam \pipeline_dffe[6] .power_up = "low";

dffeas \pipeline_dffe[7] (
	.clk(clock),
	.d(\op_1~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \pipeline_dffe[7] .is_wysiwyg = "true";
defparam \pipeline_dffe[7] .power_up = "low";

dffeas \pipeline_dffe[8] (
	.clk(clock),
	.d(\op_1~49_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \pipeline_dffe[8] .is_wysiwyg = "true";
defparam \pipeline_dffe[8] .power_up = "low";

dffeas \pipeline_dffe[9] (
	.clk(clock),
	.d(\op_1~53_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \pipeline_dffe[9] .is_wysiwyg = "true";
defparam \pipeline_dffe[9] .power_up = "low";

dffeas \pipeline_dffe[10] (
	.clk(clock),
	.d(\op_1~57_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \pipeline_dffe[10] .is_wysiwyg = "true";
defparam \pipeline_dffe[10] .power_up = "low";

dffeas \pipeline_dffe[11] (
	.clk(clock),
	.d(\op_1~61_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \pipeline_dffe[11] .is_wysiwyg = "true";
defparam \pipeline_dffe[11] .power_up = "low";

dffeas \pipeline_dffe[12] (
	.clk(clock),
	.d(\op_1~65_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_12),
	.prn(vcc));
defparam \pipeline_dffe[12] .is_wysiwyg = "true";
defparam \pipeline_dffe[12] .power_up = "low";

dffeas \pipeline_dffe[13] (
	.clk(clock),
	.d(\op_1~69_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_13),
	.prn(vcc));
defparam \pipeline_dffe[13] .is_wysiwyg = "true";
defparam \pipeline_dffe[13] .power_up = "low";

dffeas \pipeline_dffe[14] (
	.clk(clock),
	.d(\op_1~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_14),
	.prn(vcc));
defparam \pipeline_dffe[14] .is_wysiwyg = "true";
defparam \pipeline_dffe[14] .power_up = "low";

arriav_lcell_comb \op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~13_sumout ),
	.cout(\op_1~14 ),
	.shareout());
defparam \op_1~13 .extended_lut = "off";
defparam \op_1~13 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~13 .shared_arith = "off";

arriav_lcell_comb \op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_1),
	.datag(gnd),
	.cin(\op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~21_sumout ),
	.cout(\op_1~22 ),
	.shareout());
defparam \op_1~21 .extended_lut = "off";
defparam \op_1~21 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~21 .shared_arith = "off";

arriav_lcell_comb \op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_2),
	.datag(gnd),
	.cin(\op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~25_sumout ),
	.cout(\op_1~26 ),
	.shareout());
defparam \op_1~25 .extended_lut = "off";
defparam \op_1~25 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~25 .shared_arith = "off";

arriav_lcell_comb \op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~29_sumout ),
	.cout(\op_1~30 ),
	.shareout());
defparam \op_1~29 .extended_lut = "off";
defparam \op_1~29 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~29 .shared_arith = "off";

arriav_lcell_comb \op_1~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~33_sumout ),
	.cout(\op_1~34 ),
	.shareout());
defparam \op_1~33 .extended_lut = "off";
defparam \op_1~33 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~33 .shared_arith = "off";

arriav_lcell_comb \op_1~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~37_sumout ),
	.cout(\op_1~38 ),
	.shareout());
defparam \op_1~37 .extended_lut = "off";
defparam \op_1~37 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~37 .shared_arith = "off";

arriav_lcell_comb \op_1~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~41_sumout ),
	.cout(\op_1~42 ),
	.shareout());
defparam \op_1~41 .extended_lut = "off";
defparam \op_1~41 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~41 .shared_arith = "off";

arriav_lcell_comb \op_1~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~45_sumout ),
	.cout(\op_1~46 ),
	.shareout());
defparam \op_1~45 .extended_lut = "off";
defparam \op_1~45 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~45 .shared_arith = "off";

arriav_lcell_comb \op_1~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~49_sumout ),
	.cout(\op_1~50 ),
	.shareout());
defparam \op_1~49 .extended_lut = "off";
defparam \op_1~49 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~49 .shared_arith = "off";

arriav_lcell_comb \op_1~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~53_sumout ),
	.cout(\op_1~54 ),
	.shareout());
defparam \op_1~53 .extended_lut = "off";
defparam \op_1~53 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~53 .shared_arith = "off";

arriav_lcell_comb \op_1~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~57_sumout ),
	.cout(\op_1~58 ),
	.shareout());
defparam \op_1~57 .extended_lut = "off";
defparam \op_1~57 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~57 .shared_arith = "off";

arriav_lcell_comb \op_1~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~61_sumout ),
	.cout(\op_1~62 ),
	.shareout());
defparam \op_1~61 .extended_lut = "off";
defparam \op_1~61 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~61 .shared_arith = "off";

arriav_lcell_comb \op_1~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~65_sumout ),
	.cout(\op_1~66 ),
	.shareout());
defparam \op_1~65 .extended_lut = "off";
defparam \op_1~65 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~65 .shared_arith = "off";

arriav_lcell_comb \op_1~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~69_sumout ),
	.cout(\op_1~70 ),
	.shareout());
defparam \op_1~69 .extended_lut = "off";
defparam \op_1~69 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~69 .shared_arith = "off";

arriav_lcell_comb \op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~17_sumout ),
	.cout(\op_1~18 ),
	.shareout());
defparam \op_1~17 .extended_lut = "off";
defparam \op_1~17 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~17 .shared_arith = "off";

arriav_lcell_comb \op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~9_sumout ),
	.cout(\op_1~10 ),
	.shareout());
defparam \op_1~9 .extended_lut = "off";
defparam \op_1~9 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~9 .shared_arith = "off";

arriav_lcell_comb \op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_16),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~5_sumout ),
	.cout(\op_1~6 ),
	.shareout());
defparam \op_1~5 .extended_lut = "off";
defparam \op_1~5 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~5 .shared_arith = "off";

arriav_lcell_comb \op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_17),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~1_sumout ),
	.cout(),
	.shareout());
defparam \op_1~1 .extended_lut = "off";
defparam \op_1~1 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~1 .shared_arith = "off";

endmodule

module nco_test_cordic_axor_1p_lpm_12 (
	sin_o_0,
	pipeline_dffe_17,
	pipeline_dffe_16,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	pipeline_dffe_15,
	dffe16,
	dffe18,
	pipeline_dffe_171,
	dffe161,
	dffe17,
	pipeline_dffe_161,
	pipeline_dffe_151,
	pipeline_dffe_01,
	pipeline_dffe_18,
	pipeline_dffe_21,
	pipeline_dffe_31,
	pipeline_dffe_41,
	pipeline_dffe_51,
	pipeline_dffe_61,
	pipeline_dffe_71,
	pipeline_dffe_81,
	pipeline_dffe_91,
	pipeline_dffe_101,
	pipeline_dffe_111,
	pipeline_dffe_121,
	pipeline_dffe_131,
	pipeline_dffe_141,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	sin_o_0;
output 	pipeline_dffe_17;
output 	pipeline_dffe_16;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
output 	pipeline_dffe_15;
input 	dffe16;
input 	dffe18;
input 	pipeline_dffe_171;
input 	dffe161;
input 	dffe17;
input 	pipeline_dffe_161;
input 	pipeline_dffe_151;
input 	pipeline_dffe_01;
input 	pipeline_dffe_18;
input 	pipeline_dffe_21;
input 	pipeline_dffe_31;
input 	pipeline_dffe_41;
input 	pipeline_dffe_51;
input 	pipeline_dffe_61;
input 	pipeline_dffe_71;
input 	pipeline_dffe_81;
input 	pipeline_dffe_91;
input 	pipeline_dffe_101;
input 	pipeline_dffe_111;
input 	pipeline_dffe_121;
input 	pipeline_dffe_131;
input 	pipeline_dffe_141;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[17]~q ;
wire \xordvalue[10]~q ;
wire \Add0~1_sumout ;
wire \a[16]~q ;
wire \a[0]~q ;
wire \xordvalue[0]~q ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \a[15]~q ;
wire \a[1]~q ;
wire \xordvalue[1]~q ;
wire \a[2]~q ;
wire \a[3]~q ;
wire \a[4]~q ;
wire \a[5]~q ;
wire \a[6]~q ;
wire \a[7]~q ;
wire \a[8]~q ;
wire \a[9]~q ;
wire \a[10]~q ;
wire \a[11]~q ;
wire \a[12]~q ;
wire \a[13]~q ;
wire \a[14]~q ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~65_sumout ;
wire \Add0~66 ;
wire \Add0~69_sumout ;
wire \Add0~70 ;
wire \xordvalue~0_combout ;
wire \xordvalue~1_combout ;
wire \xordvalue~2_combout ;


nco_test_lpm_add_sub_14 u0(
	.a_17(\a[17]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.a_16(\a[16]~q ),
	.a_0(\a[0]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_15(\a[15]~q ),
	.a_1(\a[1]~q ),
	.xordvalue_1(\xordvalue[1]~q ),
	.a_2(\a[2]~q ),
	.a_3(\a[3]~q ),
	.a_4(\a[4]~q ),
	.a_5(\a[5]~q ),
	.a_6(\a[6]~q ),
	.a_7(\a[7]~q ),
	.a_8(\a[8]~q ),
	.a_9(\a[9]~q ),
	.a_10(\a[10]~q ),
	.a_11(\a[11]~q ),
	.a_12(\a[12]~q ),
	.a_13(\a[13]~q ),
	.a_14(\a[14]~q ),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_15(pipeline_dffe_15),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[17] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[17]~q ),
	.prn(vcc));
defparam \a[17] .is_wysiwyg = "true";
defparam \a[17] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_171),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h00000000000000FF;
defparam \Add0~1 .shared_arith = "off";

dffeas \a[16] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[16]~q ),
	.prn(vcc));
defparam \a[16] .is_wysiwyg = "true";
defparam \a[16] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h00000000000000FF;
defparam \Add0~5 .shared_arith = "off";

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \xordvalue[1] (
	.clk(clk),
	.d(\xordvalue~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[1]~q ),
	.prn(vcc));
defparam \xordvalue[1] .is_wysiwyg = "true";
defparam \xordvalue[1] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe16),
	.datae(gnd),
	.dataf(!pipeline_dffe_01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~9 .shared_arith = "off";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h00000000000000FF;
defparam \Add0~13 .shared_arith = "off";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_18),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h00000000000000FF;
defparam \Add0~17 .shared_arith = "off";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h00000000000000FF;
defparam \Add0~21 .shared_arith = "off";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h00000000000000FF;
defparam \Add0~25 .shared_arith = "off";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h00000000000000FF;
defparam \Add0~29 .shared_arith = "off";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h00000000000000FF;
defparam \Add0~33 .shared_arith = "off";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h00000000000000FF;
defparam \Add0~37 .shared_arith = "off";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h00000000000000FF;
defparam \Add0~41 .shared_arith = "off";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h00000000000000FF;
defparam \Add0~45 .shared_arith = "off";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout());
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h00000000000000FF;
defparam \Add0~49 .shared_arith = "off";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout());
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h00000000000000FF;
defparam \Add0~53 .shared_arith = "off";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout());
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h00000000000000FF;
defparam \Add0~57 .shared_arith = "off";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout());
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h00000000000000FF;
defparam \Add0~61 .shared_arith = "off";

arriav_lcell_comb \Add0~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~65_sumout ),
	.cout(\Add0~66 ),
	.shareout());
defparam \Add0~65 .extended_lut = "off";
defparam \Add0~65 .lut_mask = 64'h00000000000000FF;
defparam \Add0~65 .shared_arith = "off";

arriav_lcell_comb \Add0~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~69_sumout ),
	.cout(\Add0~70 ),
	.shareout());
defparam \Add0~69 .extended_lut = "off";
defparam \Add0~69 .lut_mask = 64'h00000000000000FF;
defparam \Add0~69 .shared_arith = "off";

arriav_lcell_comb \xordvalue~0 (
	.dataa(!dffe16),
	.datab(!dffe18),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

arriav_lcell_comb \xordvalue~1 (
	.dataa(!dffe16),
	.datab(!dffe161),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~1 .extended_lut = "off";
defparam \xordvalue~1 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~1 .shared_arith = "off";

arriav_lcell_comb \xordvalue~2 (
	.dataa(!dffe16),
	.datab(!dffe17),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~2 .extended_lut = "off";
defparam \xordvalue~2 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~2 .shared_arith = "off";

endmodule

module nco_test_lpm_add_sub_14 (
	a_17,
	xordvalue_10,
	a_16,
	a_0,
	xordvalue_0,
	a_15,
	a_1,
	xordvalue_1,
	a_2,
	a_3,
	a_4,
	a_5,
	a_6,
	a_7,
	a_8,
	a_9,
	a_10,
	a_11,
	a_12,
	a_13,
	a_14,
	pipeline_dffe_17,
	pipeline_dffe_16,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	pipeline_dffe_15,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_10;
input 	a_16;
input 	a_0;
input 	xordvalue_0;
input 	a_15;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	a_3;
input 	a_4;
input 	a_5;
input 	a_6;
input 	a_7;
input 	a_8;
input 	a_9;
input 	a_10;
input 	a_11;
input 	a_12;
input 	a_13;
input 	a_14;
output 	pipeline_dffe_17;
output 	pipeline_dffe_16;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
output 	pipeline_dffe_15;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_add_sub_0qg_12 auto_generated(
	.a_17(a_17),
	.xordvalue_10(xordvalue_10),
	.a_16(a_16),
	.a_0(a_0),
	.xordvalue_0(xordvalue_0),
	.a_15(a_15),
	.a_1(a_1),
	.xordvalue_1(xordvalue_1),
	.a_2(a_2),
	.a_3(a_3),
	.a_4(a_4),
	.a_5(a_5),
	.a_6(a_6),
	.a_7(a_7),
	.a_8(a_8),
	.a_9(a_9),
	.a_10(a_10),
	.a_11(a_11),
	.a_12(a_12),
	.a_13(a_13),
	.a_14(a_14),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_15(pipeline_dffe_15),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module nco_test_add_sub_0qg_12 (
	a_17,
	xordvalue_10,
	a_16,
	a_0,
	xordvalue_0,
	a_15,
	a_1,
	xordvalue_1,
	a_2,
	a_3,
	a_4,
	a_5,
	a_6,
	a_7,
	a_8,
	a_9,
	a_10,
	a_11,
	a_12,
	a_13,
	a_14,
	pipeline_dffe_17,
	pipeline_dffe_16,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	pipeline_dffe_15,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_10;
input 	a_16;
input 	a_0;
input 	xordvalue_0;
input 	a_15;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	a_3;
input 	a_4;
input 	a_5;
input 	a_6;
input 	a_7;
input 	a_8;
input 	a_9;
input 	a_10;
input 	a_11;
input 	a_12;
input 	a_13;
input 	a_14;
output 	pipeline_dffe_17;
output 	pipeline_dffe_16;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
output 	pipeline_dffe_15;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \op_1~10 ;
wire \op_1~18 ;
wire \op_1~22 ;
wire \op_1~26 ;
wire \op_1~30 ;
wire \op_1~34 ;
wire \op_1~38 ;
wire \op_1~42 ;
wire \op_1~46 ;
wire \op_1~50 ;
wire \op_1~54 ;
wire \op_1~58 ;
wire \op_1~62 ;
wire \op_1~66 ;
wire \op_1~70 ;
wire \op_1~14 ;
wire \op_1~6 ;
wire \op_1~1_sumout ;
wire \op_1~5_sumout ;
wire \op_1~9_sumout ;
wire \op_1~17_sumout ;
wire \op_1~21_sumout ;
wire \op_1~25_sumout ;
wire \op_1~29_sumout ;
wire \op_1~33_sumout ;
wire \op_1~37_sumout ;
wire \op_1~41_sumout ;
wire \op_1~45_sumout ;
wire \op_1~49_sumout ;
wire \op_1~53_sumout ;
wire \op_1~57_sumout ;
wire \op_1~61_sumout ;
wire \op_1~65_sumout ;
wire \op_1~69_sumout ;
wire \op_1~13_sumout ;


dffeas \pipeline_dffe[17] (
	.clk(clock),
	.d(\op_1~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_17),
	.prn(vcc));
defparam \pipeline_dffe[17] .is_wysiwyg = "true";
defparam \pipeline_dffe[17] .power_up = "low";

dffeas \pipeline_dffe[16] (
	.clk(clock),
	.d(\op_1~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_16),
	.prn(vcc));
defparam \pipeline_dffe[16] .is_wysiwyg = "true";
defparam \pipeline_dffe[16] .power_up = "low";

dffeas \pipeline_dffe[0] (
	.clk(clock),
	.d(\op_1~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_0),
	.prn(vcc));
defparam \pipeline_dffe[0] .is_wysiwyg = "true";
defparam \pipeline_dffe[0] .power_up = "low";

dffeas \pipeline_dffe[1] (
	.clk(clock),
	.d(\op_1~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_1),
	.prn(vcc));
defparam \pipeline_dffe[1] .is_wysiwyg = "true";
defparam \pipeline_dffe[1] .power_up = "low";

dffeas \pipeline_dffe[2] (
	.clk(clock),
	.d(\op_1~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \pipeline_dffe[2] .is_wysiwyg = "true";
defparam \pipeline_dffe[2] .power_up = "low";

dffeas \pipeline_dffe[3] (
	.clk(clock),
	.d(\op_1~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \pipeline_dffe[3] .is_wysiwyg = "true";
defparam \pipeline_dffe[3] .power_up = "low";

dffeas \pipeline_dffe[4] (
	.clk(clock),
	.d(\op_1~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \pipeline_dffe[4] .is_wysiwyg = "true";
defparam \pipeline_dffe[4] .power_up = "low";

dffeas \pipeline_dffe[5] (
	.clk(clock),
	.d(\op_1~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \pipeline_dffe[5] .is_wysiwyg = "true";
defparam \pipeline_dffe[5] .power_up = "low";

dffeas \pipeline_dffe[6] (
	.clk(clock),
	.d(\op_1~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \pipeline_dffe[6] .is_wysiwyg = "true";
defparam \pipeline_dffe[6] .power_up = "low";

dffeas \pipeline_dffe[7] (
	.clk(clock),
	.d(\op_1~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \pipeline_dffe[7] .is_wysiwyg = "true";
defparam \pipeline_dffe[7] .power_up = "low";

dffeas \pipeline_dffe[8] (
	.clk(clock),
	.d(\op_1~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \pipeline_dffe[8] .is_wysiwyg = "true";
defparam \pipeline_dffe[8] .power_up = "low";

dffeas \pipeline_dffe[9] (
	.clk(clock),
	.d(\op_1~49_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \pipeline_dffe[9] .is_wysiwyg = "true";
defparam \pipeline_dffe[9] .power_up = "low";

dffeas \pipeline_dffe[10] (
	.clk(clock),
	.d(\op_1~53_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \pipeline_dffe[10] .is_wysiwyg = "true";
defparam \pipeline_dffe[10] .power_up = "low";

dffeas \pipeline_dffe[11] (
	.clk(clock),
	.d(\op_1~57_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \pipeline_dffe[11] .is_wysiwyg = "true";
defparam \pipeline_dffe[11] .power_up = "low";

dffeas \pipeline_dffe[12] (
	.clk(clock),
	.d(\op_1~61_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_12),
	.prn(vcc));
defparam \pipeline_dffe[12] .is_wysiwyg = "true";
defparam \pipeline_dffe[12] .power_up = "low";

dffeas \pipeline_dffe[13] (
	.clk(clock),
	.d(\op_1~65_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_13),
	.prn(vcc));
defparam \pipeline_dffe[13] .is_wysiwyg = "true";
defparam \pipeline_dffe[13] .power_up = "low";

dffeas \pipeline_dffe[14] (
	.clk(clock),
	.d(\op_1~69_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_14),
	.prn(vcc));
defparam \pipeline_dffe[14] .is_wysiwyg = "true";
defparam \pipeline_dffe[14] .power_up = "low";

dffeas \pipeline_dffe[15] (
	.clk(clock),
	.d(\op_1~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_15),
	.prn(vcc));
defparam \pipeline_dffe[15] .is_wysiwyg = "true";
defparam \pipeline_dffe[15] .power_up = "low";

arriav_lcell_comb \op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~9_sumout ),
	.cout(\op_1~10 ),
	.shareout());
defparam \op_1~9 .extended_lut = "off";
defparam \op_1~9 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~9 .shared_arith = "off";

arriav_lcell_comb \op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_1),
	.datag(gnd),
	.cin(\op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~17_sumout ),
	.cout(\op_1~18 ),
	.shareout());
defparam \op_1~17 .extended_lut = "off";
defparam \op_1~17 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~17 .shared_arith = "off";

arriav_lcell_comb \op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~21_sumout ),
	.cout(\op_1~22 ),
	.shareout());
defparam \op_1~21 .extended_lut = "off";
defparam \op_1~21 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~21 .shared_arith = "off";

arriav_lcell_comb \op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~25_sumout ),
	.cout(\op_1~26 ),
	.shareout());
defparam \op_1~25 .extended_lut = "off";
defparam \op_1~25 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~25 .shared_arith = "off";

arriav_lcell_comb \op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~29_sumout ),
	.cout(\op_1~30 ),
	.shareout());
defparam \op_1~29 .extended_lut = "off";
defparam \op_1~29 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~29 .shared_arith = "off";

arriav_lcell_comb \op_1~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~33_sumout ),
	.cout(\op_1~34 ),
	.shareout());
defparam \op_1~33 .extended_lut = "off";
defparam \op_1~33 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~33 .shared_arith = "off";

arriav_lcell_comb \op_1~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~37_sumout ),
	.cout(\op_1~38 ),
	.shareout());
defparam \op_1~37 .extended_lut = "off";
defparam \op_1~37 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~37 .shared_arith = "off";

arriav_lcell_comb \op_1~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~41_sumout ),
	.cout(\op_1~42 ),
	.shareout());
defparam \op_1~41 .extended_lut = "off";
defparam \op_1~41 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~41 .shared_arith = "off";

arriav_lcell_comb \op_1~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~45_sumout ),
	.cout(\op_1~46 ),
	.shareout());
defparam \op_1~45 .extended_lut = "off";
defparam \op_1~45 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~45 .shared_arith = "off";

arriav_lcell_comb \op_1~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~49_sumout ),
	.cout(\op_1~50 ),
	.shareout());
defparam \op_1~49 .extended_lut = "off";
defparam \op_1~49 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~49 .shared_arith = "off";

arriav_lcell_comb \op_1~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~53_sumout ),
	.cout(\op_1~54 ),
	.shareout());
defparam \op_1~53 .extended_lut = "off";
defparam \op_1~53 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~53 .shared_arith = "off";

arriav_lcell_comb \op_1~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~57_sumout ),
	.cout(\op_1~58 ),
	.shareout());
defparam \op_1~57 .extended_lut = "off";
defparam \op_1~57 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~57 .shared_arith = "off";

arriav_lcell_comb \op_1~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~61_sumout ),
	.cout(\op_1~62 ),
	.shareout());
defparam \op_1~61 .extended_lut = "off";
defparam \op_1~61 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~61 .shared_arith = "off";

arriav_lcell_comb \op_1~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~65_sumout ),
	.cout(\op_1~66 ),
	.shareout());
defparam \op_1~65 .extended_lut = "off";
defparam \op_1~65 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~65 .shared_arith = "off";

arriav_lcell_comb \op_1~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~69_sumout ),
	.cout(\op_1~70 ),
	.shareout());
defparam \op_1~69 .extended_lut = "off";
defparam \op_1~69 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~69 .shared_arith = "off";

arriav_lcell_comb \op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~13_sumout ),
	.cout(\op_1~14 ),
	.shareout());
defparam \op_1~13 .extended_lut = "off";
defparam \op_1~13 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~13 .shared_arith = "off";

arriav_lcell_comb \op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_16),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~5_sumout ),
	.cout(\op_1~6 ),
	.shareout());
defparam \op_1~5 .extended_lut = "off";
defparam \op_1~5 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~5 .shared_arith = "off";

arriav_lcell_comb \op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_17),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~1_sumout ),
	.cout(),
	.shareout());
defparam \op_1~1 .extended_lut = "off";
defparam \op_1~1 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~1 .shared_arith = "off";

endmodule

module nco_test_cordic_axor_1p_lpm_13 (
	a_0,
	xordvalue_11,
	cor1x_10,
	sin_o_0,
	pipeline_dffe_17,
	pipeline_dffe_16,
	dffe16,
	xordvalue,
	pipeline_dffe_15,
	pipeline_dffe_14,
	pipeline_dffe_13,
	pipeline_dffe_12,
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_7,
	pipeline_dffe_6,
	pipeline_dffe_5,
	pipeline_dffe_4,
	pipeline_dffe_3,
	pipeline_dffe_2,
	pipeline_dffe_1,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	a_0;
output 	xordvalue_11;
input 	cor1x_10;
input 	sin_o_0;
output 	pipeline_dffe_17;
output 	pipeline_dffe_16;
input 	dffe16;
output 	xordvalue;
output 	pipeline_dffe_15;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_7;
output 	pipeline_dffe_6;
output 	pipeline_dffe_5;
output 	pipeline_dffe_4;
output 	pipeline_dffe_3;
output 	pipeline_dffe_2;
output 	pipeline_dffe_1;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[10]~q ;


nco_test_lpm_add_sub_17 u0(
	.a_0(a_0),
	.xordvalue_11(xordvalue_11),
	.a_10(\a[10]~q ),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_1(pipeline_dffe_1),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[10] (
	.clk(clk),
	.d(cor1x_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(dffe16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(a_0),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \xordvalue[11] (
	.clk(clk),
	.d(xordvalue),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(xordvalue_11),
	.prn(vcc));
defparam \xordvalue[11] .is_wysiwyg = "true";
defparam \xordvalue[11] .power_up = "low";

arriav_lcell_comb \xordvalue~0 (
	.dataa(!dffe16),
	.datab(!cor1x_10),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(xordvalue),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

endmodule

module nco_test_cordic_axor_1p_lpm_14 (
	sin_o_0,
	pipeline_dffe_17,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	pipeline_dffe_15,
	pipeline_dffe_16,
	dffe16,
	pipeline_dffe_171,
	dffe18,
	dffe17,
	pipeline_dffe_161,
	pipeline_dffe_01,
	pipeline_dffe_18,
	pipeline_dffe_21,
	pipeline_dffe_31,
	pipeline_dffe_41,
	pipeline_dffe_51,
	pipeline_dffe_61,
	pipeline_dffe_71,
	pipeline_dffe_81,
	pipeline_dffe_91,
	pipeline_dffe_101,
	pipeline_dffe_111,
	pipeline_dffe_121,
	pipeline_dffe_131,
	pipeline_dffe_141,
	pipeline_dffe_151,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	sin_o_0;
output 	pipeline_dffe_17;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
output 	pipeline_dffe_15;
output 	pipeline_dffe_16;
input 	dffe16;
input 	pipeline_dffe_171;
input 	dffe18;
input 	dffe17;
input 	pipeline_dffe_161;
input 	pipeline_dffe_01;
input 	pipeline_dffe_18;
input 	pipeline_dffe_21;
input 	pipeline_dffe_31;
input 	pipeline_dffe_41;
input 	pipeline_dffe_51;
input 	pipeline_dffe_61;
input 	pipeline_dffe_71;
input 	pipeline_dffe_81;
input 	pipeline_dffe_91;
input 	pipeline_dffe_101;
input 	pipeline_dffe_111;
input 	pipeline_dffe_121;
input 	pipeline_dffe_131;
input 	pipeline_dffe_141;
input 	pipeline_dffe_151;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[17]~q ;
wire \xordvalue[10]~q ;
wire \a[0]~q ;
wire \xordvalue[0]~q ;
wire \Add0~1_sumout ;
wire \a[16]~q ;
wire \a[1]~q ;
wire \a[2]~q ;
wire \a[3]~q ;
wire \a[4]~q ;
wire \a[5]~q ;
wire \a[6]~q ;
wire \a[7]~q ;
wire \a[8]~q ;
wire \a[9]~q ;
wire \a[10]~q ;
wire \a[11]~q ;
wire \a[12]~q ;
wire \a[13]~q ;
wire \a[14]~q ;
wire \a[15]~q ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~65_sumout ;
wire \Add0~66 ;
wire \Add0~69_sumout ;
wire \Add0~70 ;
wire \xordvalue~0_combout ;
wire \xordvalue~1_combout ;


nco_test_lpm_add_sub_15 u0(
	.a_17(\a[17]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.a_0(\a[0]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_16(\a[16]~q ),
	.a_1(\a[1]~q ),
	.a_2(\a[2]~q ),
	.a_3(\a[3]~q ),
	.a_4(\a[4]~q ),
	.a_5(\a[5]~q ),
	.a_6(\a[6]~q ),
	.a_7(\a[7]~q ),
	.a_8(\a[8]~q ),
	.a_9(\a[9]~q ),
	.a_10(\a[10]~q ),
	.a_11(\a[11]~q ),
	.a_12(\a[12]~q ),
	.a_13(\a[13]~q ),
	.a_14(\a[14]~q ),
	.a_15(\a[15]~q ),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_16(pipeline_dffe_16),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[17] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[17]~q ),
	.prn(vcc));
defparam \a[17] .is_wysiwyg = "true";
defparam \a[17] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_171),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h00000000000000FF;
defparam \Add0~1 .shared_arith = "off";

dffeas \a[16] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[16]~q ),
	.prn(vcc));
defparam \a[16] .is_wysiwyg = "true";
defparam \a[16] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe16),
	.datae(gnd),
	.dataf(!pipeline_dffe_01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~5 .shared_arith = "off";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h00000000000000FF;
defparam \Add0~9 .shared_arith = "off";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_18),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h00000000000000FF;
defparam \Add0~13 .shared_arith = "off";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h00000000000000FF;
defparam \Add0~17 .shared_arith = "off";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h00000000000000FF;
defparam \Add0~21 .shared_arith = "off";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h00000000000000FF;
defparam \Add0~25 .shared_arith = "off";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h00000000000000FF;
defparam \Add0~29 .shared_arith = "off";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h00000000000000FF;
defparam \Add0~33 .shared_arith = "off";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h00000000000000FF;
defparam \Add0~37 .shared_arith = "off";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h00000000000000FF;
defparam \Add0~41 .shared_arith = "off";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h00000000000000FF;
defparam \Add0~45 .shared_arith = "off";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout());
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h00000000000000FF;
defparam \Add0~49 .shared_arith = "off";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout());
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h00000000000000FF;
defparam \Add0~53 .shared_arith = "off";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout());
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h00000000000000FF;
defparam \Add0~57 .shared_arith = "off";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout());
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h00000000000000FF;
defparam \Add0~61 .shared_arith = "off";

arriav_lcell_comb \Add0~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~65_sumout ),
	.cout(\Add0~66 ),
	.shareout());
defparam \Add0~65 .extended_lut = "off";
defparam \Add0~65 .lut_mask = 64'h00000000000000FF;
defparam \Add0~65 .shared_arith = "off";

arriav_lcell_comb \Add0~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~69_sumout ),
	.cout(\Add0~70 ),
	.shareout());
defparam \Add0~69 .extended_lut = "off";
defparam \Add0~69 .lut_mask = 64'h00000000000000FF;
defparam \Add0~69 .shared_arith = "off";

arriav_lcell_comb \xordvalue~0 (
	.dataa(!dffe18),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

arriav_lcell_comb \xordvalue~1 (
	.dataa(!dffe17),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~1 .extended_lut = "off";
defparam \xordvalue~1 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~1 .shared_arith = "off";

endmodule

module nco_test_lpm_add_sub_15 (
	a_17,
	xordvalue_10,
	a_0,
	xordvalue_0,
	a_16,
	a_1,
	a_2,
	a_3,
	a_4,
	a_5,
	a_6,
	a_7,
	a_8,
	a_9,
	a_10,
	a_11,
	a_12,
	a_13,
	a_14,
	a_15,
	pipeline_dffe_17,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	pipeline_dffe_15,
	pipeline_dffe_16,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_10;
input 	a_0;
input 	xordvalue_0;
input 	a_16;
input 	a_1;
input 	a_2;
input 	a_3;
input 	a_4;
input 	a_5;
input 	a_6;
input 	a_7;
input 	a_8;
input 	a_9;
input 	a_10;
input 	a_11;
input 	a_12;
input 	a_13;
input 	a_14;
input 	a_15;
output 	pipeline_dffe_17;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
output 	pipeline_dffe_15;
output 	pipeline_dffe_16;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_add_sub_0qg_13 auto_generated(
	.a_17(a_17),
	.xordvalue_10(xordvalue_10),
	.a_0(a_0),
	.xordvalue_0(xordvalue_0),
	.a_16(a_16),
	.a_1(a_1),
	.a_2(a_2),
	.a_3(a_3),
	.a_4(a_4),
	.a_5(a_5),
	.a_6(a_6),
	.a_7(a_7),
	.a_8(a_8),
	.a_9(a_9),
	.a_10(a_10),
	.a_11(a_11),
	.a_12(a_12),
	.a_13(a_13),
	.a_14(a_14),
	.a_15(a_15),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_16(pipeline_dffe_16),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module nco_test_add_sub_0qg_13 (
	a_17,
	xordvalue_10,
	a_0,
	xordvalue_0,
	a_16,
	a_1,
	a_2,
	a_3,
	a_4,
	a_5,
	a_6,
	a_7,
	a_8,
	a_9,
	a_10,
	a_11,
	a_12,
	a_13,
	a_14,
	a_15,
	pipeline_dffe_17,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	pipeline_dffe_15,
	pipeline_dffe_16,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_10;
input 	a_0;
input 	xordvalue_0;
input 	a_16;
input 	a_1;
input 	a_2;
input 	a_3;
input 	a_4;
input 	a_5;
input 	a_6;
input 	a_7;
input 	a_8;
input 	a_9;
input 	a_10;
input 	a_11;
input 	a_12;
input 	a_13;
input 	a_14;
input 	a_15;
output 	pipeline_dffe_17;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
output 	pipeline_dffe_15;
output 	pipeline_dffe_16;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \op_1~6 ;
wire \op_1~14 ;
wire \op_1~18 ;
wire \op_1~22 ;
wire \op_1~26 ;
wire \op_1~30 ;
wire \op_1~34 ;
wire \op_1~38 ;
wire \op_1~42 ;
wire \op_1~46 ;
wire \op_1~50 ;
wire \op_1~54 ;
wire \op_1~58 ;
wire \op_1~62 ;
wire \op_1~66 ;
wire \op_1~70 ;
wire \op_1~10 ;
wire \op_1~1_sumout ;
wire \op_1~5_sumout ;
wire \op_1~13_sumout ;
wire \op_1~17_sumout ;
wire \op_1~21_sumout ;
wire \op_1~25_sumout ;
wire \op_1~29_sumout ;
wire \op_1~33_sumout ;
wire \op_1~37_sumout ;
wire \op_1~41_sumout ;
wire \op_1~45_sumout ;
wire \op_1~49_sumout ;
wire \op_1~53_sumout ;
wire \op_1~57_sumout ;
wire \op_1~61_sumout ;
wire \op_1~65_sumout ;
wire \op_1~69_sumout ;
wire \op_1~9_sumout ;


dffeas \pipeline_dffe[17] (
	.clk(clock),
	.d(\op_1~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_17),
	.prn(vcc));
defparam \pipeline_dffe[17] .is_wysiwyg = "true";
defparam \pipeline_dffe[17] .power_up = "low";

dffeas \pipeline_dffe[0] (
	.clk(clock),
	.d(\op_1~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_0),
	.prn(vcc));
defparam \pipeline_dffe[0] .is_wysiwyg = "true";
defparam \pipeline_dffe[0] .power_up = "low";

dffeas \pipeline_dffe[1] (
	.clk(clock),
	.d(\op_1~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_1),
	.prn(vcc));
defparam \pipeline_dffe[1] .is_wysiwyg = "true";
defparam \pipeline_dffe[1] .power_up = "low";

dffeas \pipeline_dffe[2] (
	.clk(clock),
	.d(\op_1~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \pipeline_dffe[2] .is_wysiwyg = "true";
defparam \pipeline_dffe[2] .power_up = "low";

dffeas \pipeline_dffe[3] (
	.clk(clock),
	.d(\op_1~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \pipeline_dffe[3] .is_wysiwyg = "true";
defparam \pipeline_dffe[3] .power_up = "low";

dffeas \pipeline_dffe[4] (
	.clk(clock),
	.d(\op_1~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \pipeline_dffe[4] .is_wysiwyg = "true";
defparam \pipeline_dffe[4] .power_up = "low";

dffeas \pipeline_dffe[5] (
	.clk(clock),
	.d(\op_1~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \pipeline_dffe[5] .is_wysiwyg = "true";
defparam \pipeline_dffe[5] .power_up = "low";

dffeas \pipeline_dffe[6] (
	.clk(clock),
	.d(\op_1~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \pipeline_dffe[6] .is_wysiwyg = "true";
defparam \pipeline_dffe[6] .power_up = "low";

dffeas \pipeline_dffe[7] (
	.clk(clock),
	.d(\op_1~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \pipeline_dffe[7] .is_wysiwyg = "true";
defparam \pipeline_dffe[7] .power_up = "low";

dffeas \pipeline_dffe[8] (
	.clk(clock),
	.d(\op_1~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \pipeline_dffe[8] .is_wysiwyg = "true";
defparam \pipeline_dffe[8] .power_up = "low";

dffeas \pipeline_dffe[9] (
	.clk(clock),
	.d(\op_1~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \pipeline_dffe[9] .is_wysiwyg = "true";
defparam \pipeline_dffe[9] .power_up = "low";

dffeas \pipeline_dffe[10] (
	.clk(clock),
	.d(\op_1~49_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \pipeline_dffe[10] .is_wysiwyg = "true";
defparam \pipeline_dffe[10] .power_up = "low";

dffeas \pipeline_dffe[11] (
	.clk(clock),
	.d(\op_1~53_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \pipeline_dffe[11] .is_wysiwyg = "true";
defparam \pipeline_dffe[11] .power_up = "low";

dffeas \pipeline_dffe[12] (
	.clk(clock),
	.d(\op_1~57_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_12),
	.prn(vcc));
defparam \pipeline_dffe[12] .is_wysiwyg = "true";
defparam \pipeline_dffe[12] .power_up = "low";

dffeas \pipeline_dffe[13] (
	.clk(clock),
	.d(\op_1~61_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_13),
	.prn(vcc));
defparam \pipeline_dffe[13] .is_wysiwyg = "true";
defparam \pipeline_dffe[13] .power_up = "low";

dffeas \pipeline_dffe[14] (
	.clk(clock),
	.d(\op_1~65_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_14),
	.prn(vcc));
defparam \pipeline_dffe[14] .is_wysiwyg = "true";
defparam \pipeline_dffe[14] .power_up = "low";

dffeas \pipeline_dffe[15] (
	.clk(clock),
	.d(\op_1~69_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_15),
	.prn(vcc));
defparam \pipeline_dffe[15] .is_wysiwyg = "true";
defparam \pipeline_dffe[15] .power_up = "low";

dffeas \pipeline_dffe[16] (
	.clk(clock),
	.d(\op_1~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_16),
	.prn(vcc));
defparam \pipeline_dffe[16] .is_wysiwyg = "true";
defparam \pipeline_dffe[16] .power_up = "low";

arriav_lcell_comb \op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~5_sumout ),
	.cout(\op_1~6 ),
	.shareout());
defparam \op_1~5 .extended_lut = "off";
defparam \op_1~5 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~5 .shared_arith = "off";

arriav_lcell_comb \op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~13_sumout ),
	.cout(\op_1~14 ),
	.shareout());
defparam \op_1~13 .extended_lut = "off";
defparam \op_1~13 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~13 .shared_arith = "off";

arriav_lcell_comb \op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~17_sumout ),
	.cout(\op_1~18 ),
	.shareout());
defparam \op_1~17 .extended_lut = "off";
defparam \op_1~17 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~17 .shared_arith = "off";

arriav_lcell_comb \op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~21_sumout ),
	.cout(\op_1~22 ),
	.shareout());
defparam \op_1~21 .extended_lut = "off";
defparam \op_1~21 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~21 .shared_arith = "off";

arriav_lcell_comb \op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~25_sumout ),
	.cout(\op_1~26 ),
	.shareout());
defparam \op_1~25 .extended_lut = "off";
defparam \op_1~25 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~25 .shared_arith = "off";

arriav_lcell_comb \op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~29_sumout ),
	.cout(\op_1~30 ),
	.shareout());
defparam \op_1~29 .extended_lut = "off";
defparam \op_1~29 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~29 .shared_arith = "off";

arriav_lcell_comb \op_1~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~33_sumout ),
	.cout(\op_1~34 ),
	.shareout());
defparam \op_1~33 .extended_lut = "off";
defparam \op_1~33 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~33 .shared_arith = "off";

arriav_lcell_comb \op_1~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~37_sumout ),
	.cout(\op_1~38 ),
	.shareout());
defparam \op_1~37 .extended_lut = "off";
defparam \op_1~37 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~37 .shared_arith = "off";

arriav_lcell_comb \op_1~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~41_sumout ),
	.cout(\op_1~42 ),
	.shareout());
defparam \op_1~41 .extended_lut = "off";
defparam \op_1~41 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~41 .shared_arith = "off";

arriav_lcell_comb \op_1~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~45_sumout ),
	.cout(\op_1~46 ),
	.shareout());
defparam \op_1~45 .extended_lut = "off";
defparam \op_1~45 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~45 .shared_arith = "off";

arriav_lcell_comb \op_1~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~49_sumout ),
	.cout(\op_1~50 ),
	.shareout());
defparam \op_1~49 .extended_lut = "off";
defparam \op_1~49 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~49 .shared_arith = "off";

arriav_lcell_comb \op_1~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~53_sumout ),
	.cout(\op_1~54 ),
	.shareout());
defparam \op_1~53 .extended_lut = "off";
defparam \op_1~53 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~53 .shared_arith = "off";

arriav_lcell_comb \op_1~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~57_sumout ),
	.cout(\op_1~58 ),
	.shareout());
defparam \op_1~57 .extended_lut = "off";
defparam \op_1~57 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~57 .shared_arith = "off";

arriav_lcell_comb \op_1~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~61_sumout ),
	.cout(\op_1~62 ),
	.shareout());
defparam \op_1~61 .extended_lut = "off";
defparam \op_1~61 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~61 .shared_arith = "off";

arriav_lcell_comb \op_1~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~65_sumout ),
	.cout(\op_1~66 ),
	.shareout());
defparam \op_1~65 .extended_lut = "off";
defparam \op_1~65 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~65 .shared_arith = "off";

arriav_lcell_comb \op_1~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~69_sumout ),
	.cout(\op_1~70 ),
	.shareout());
defparam \op_1~69 .extended_lut = "off";
defparam \op_1~69 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~69 .shared_arith = "off";

arriav_lcell_comb \op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_16),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~9_sumout ),
	.cout(\op_1~10 ),
	.shareout());
defparam \op_1~9 .extended_lut = "off";
defparam \op_1~9 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~9 .shared_arith = "off";

arriav_lcell_comb \op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_17),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~1_sumout ),
	.cout(),
	.shareout());
defparam \op_1~1 .extended_lut = "off";
defparam \op_1~1 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~1 .shared_arith = "off";

endmodule

module nco_test_cordic_axor_1p_lpm_15 (
	sin_o_0,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	pipeline_dffe_15,
	pipeline_dffe_16,
	pipeline_dffe_17,
	dffe16,
	dffe18,
	pipeline_dffe_171,
	pipeline_dffe_01,
	pipeline_dffe_18,
	pipeline_dffe_21,
	pipeline_dffe_31,
	pipeline_dffe_41,
	pipeline_dffe_51,
	pipeline_dffe_61,
	pipeline_dffe_71,
	pipeline_dffe_81,
	pipeline_dffe_91,
	pipeline_dffe_101,
	pipeline_dffe_111,
	pipeline_dffe_121,
	pipeline_dffe_131,
	pipeline_dffe_141,
	pipeline_dffe_151,
	pipeline_dffe_161,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	sin_o_0;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
output 	pipeline_dffe_15;
output 	pipeline_dffe_16;
output 	pipeline_dffe_17;
input 	dffe16;
input 	dffe18;
input 	pipeline_dffe_171;
input 	pipeline_dffe_01;
input 	pipeline_dffe_18;
input 	pipeline_dffe_21;
input 	pipeline_dffe_31;
input 	pipeline_dffe_41;
input 	pipeline_dffe_51;
input 	pipeline_dffe_61;
input 	pipeline_dffe_71;
input 	pipeline_dffe_81;
input 	pipeline_dffe_91;
input 	pipeline_dffe_101;
input 	pipeline_dffe_111;
input 	pipeline_dffe_121;
input 	pipeline_dffe_131;
input 	pipeline_dffe_141;
input 	pipeline_dffe_151;
input 	pipeline_dffe_161;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[0]~q ;
wire \xordvalue[0]~q ;
wire \a[1]~q ;
wire \a[2]~q ;
wire \a[3]~q ;
wire \a[4]~q ;
wire \a[5]~q ;
wire \a[6]~q ;
wire \a[7]~q ;
wire \a[8]~q ;
wire \a[9]~q ;
wire \a[10]~q ;
wire \a[11]~q ;
wire \a[12]~q ;
wire \a[13]~q ;
wire \a[14]~q ;
wire \a[15]~q ;
wire \a[16]~q ;
wire \a[17]~q ;
wire \Add0~1_sumout ;
wire \Add0~2 ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~65_sumout ;
wire \Add0~66 ;
wire \Add0~69_sumout ;
wire \xordvalue~0_combout ;


nco_test_lpm_add_sub_16 u0(
	.a_0(\a[0]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_1(\a[1]~q ),
	.a_2(\a[2]~q ),
	.a_3(\a[3]~q ),
	.a_4(\a[4]~q ),
	.a_5(\a[5]~q ),
	.a_6(\a[6]~q ),
	.a_7(\a[7]~q ),
	.a_8(\a[8]~q ),
	.a_9(\a[9]~q ),
	.a_10(\a[10]~q ),
	.a_11(\a[11]~q ),
	.a_12(\a[12]~q ),
	.a_13(\a[13]~q ),
	.a_14(\a[14]~q ),
	.a_15(\a[15]~q ),
	.a_16(\a[16]~q ),
	.a_17(\a[17]~q ),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_17(pipeline_dffe_17),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

dffeas \a[16] (
	.clk(clk),
	.d(\Add0~65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[16]~q ),
	.prn(vcc));
defparam \a[16] .is_wysiwyg = "true";
defparam \a[16] .power_up = "low";

dffeas \a[17] (
	.clk(clk),
	.d(\Add0~69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[17]~q ),
	.prn(vcc));
defparam \a[17] .is_wysiwyg = "true";
defparam \a[17] .power_up = "low";

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe16),
	.datae(gnd),
	.dataf(!pipeline_dffe_01),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF00000000FF;
defparam \Add0~1 .shared_arith = "off";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_18),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout());
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h00000000000000FF;
defparam \Add0~5 .shared_arith = "off";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout());
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h00000000000000FF;
defparam \Add0~9 .shared_arith = "off";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout());
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h00000000000000FF;
defparam \Add0~13 .shared_arith = "off";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout());
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h00000000000000FF;
defparam \Add0~17 .shared_arith = "off";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout());
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h00000000000000FF;
defparam \Add0~21 .shared_arith = "off";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout());
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h00000000000000FF;
defparam \Add0~25 .shared_arith = "off";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout());
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h00000000000000FF;
defparam \Add0~29 .shared_arith = "off";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout());
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h00000000000000FF;
defparam \Add0~33 .shared_arith = "off";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout());
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h00000000000000FF;
defparam \Add0~37 .shared_arith = "off";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout());
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h00000000000000FF;
defparam \Add0~41 .shared_arith = "off";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout());
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h00000000000000FF;
defparam \Add0~45 .shared_arith = "off";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout());
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h00000000000000FF;
defparam \Add0~49 .shared_arith = "off";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout());
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h00000000000000FF;
defparam \Add0~53 .shared_arith = "off";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout());
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h00000000000000FF;
defparam \Add0~57 .shared_arith = "off";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout());
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h00000000000000FF;
defparam \Add0~61 .shared_arith = "off";

arriav_lcell_comb \Add0~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~65_sumout ),
	.cout(\Add0~66 ),
	.shareout());
defparam \Add0~65 .extended_lut = "off";
defparam \Add0~65 .lut_mask = 64'h00000000000000FF;
defparam \Add0~65 .shared_arith = "off";

arriav_lcell_comb \Add0~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!pipeline_dffe_171),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~69_sumout ),
	.cout(),
	.shareout());
defparam \Add0~69 .extended_lut = "off";
defparam \Add0~69 .lut_mask = 64'h00000000000000FF;
defparam \Add0~69 .shared_arith = "off";

arriav_lcell_comb \xordvalue~0 (
	.dataa(!dffe16),
	.datab(!dffe18),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

endmodule

module nco_test_lpm_add_sub_16 (
	a_0,
	xordvalue_0,
	a_1,
	a_2,
	a_3,
	a_4,
	a_5,
	a_6,
	a_7,
	a_8,
	a_9,
	a_10,
	a_11,
	a_12,
	a_13,
	a_14,
	a_15,
	a_16,
	a_17,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	pipeline_dffe_15,
	pipeline_dffe_16,
	pipeline_dffe_17,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_0;
input 	xordvalue_0;
input 	a_1;
input 	a_2;
input 	a_3;
input 	a_4;
input 	a_5;
input 	a_6;
input 	a_7;
input 	a_8;
input 	a_9;
input 	a_10;
input 	a_11;
input 	a_12;
input 	a_13;
input 	a_14;
input 	a_15;
input 	a_16;
input 	a_17;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
output 	pipeline_dffe_15;
output 	pipeline_dffe_16;
output 	pipeline_dffe_17;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_add_sub_0qg_14 auto_generated(
	.a_0(a_0),
	.xordvalue_0(xordvalue_0),
	.a_1(a_1),
	.a_2(a_2),
	.a_3(a_3),
	.a_4(a_4),
	.a_5(a_5),
	.a_6(a_6),
	.a_7(a_7),
	.a_8(a_8),
	.a_9(a_9),
	.a_10(a_10),
	.a_11(a_11),
	.a_12(a_12),
	.a_13(a_13),
	.a_14(a_14),
	.a_15(a_15),
	.a_16(a_16),
	.a_17(a_17),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_17(pipeline_dffe_17),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module nco_test_add_sub_0qg_14 (
	a_0,
	xordvalue_0,
	a_1,
	a_2,
	a_3,
	a_4,
	a_5,
	a_6,
	a_7,
	a_8,
	a_9,
	a_10,
	a_11,
	a_12,
	a_13,
	a_14,
	a_15,
	a_16,
	a_17,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	pipeline_dffe_10,
	pipeline_dffe_11,
	pipeline_dffe_12,
	pipeline_dffe_13,
	pipeline_dffe_14,
	pipeline_dffe_15,
	pipeline_dffe_16,
	pipeline_dffe_17,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_0;
input 	xordvalue_0;
input 	a_1;
input 	a_2;
input 	a_3;
input 	a_4;
input 	a_5;
input 	a_6;
input 	a_7;
input 	a_8;
input 	a_9;
input 	a_10;
input 	a_11;
input 	a_12;
input 	a_13;
input 	a_14;
input 	a_15;
input 	a_16;
input 	a_17;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
output 	pipeline_dffe_10;
output 	pipeline_dffe_11;
output 	pipeline_dffe_12;
output 	pipeline_dffe_13;
output 	pipeline_dffe_14;
output 	pipeline_dffe_15;
output 	pipeline_dffe_16;
output 	pipeline_dffe_17;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \op_1~1_sumout ;
wire \op_1~2 ;
wire \op_1~5_sumout ;
wire \op_1~6 ;
wire \op_1~9_sumout ;
wire \op_1~10 ;
wire \op_1~13_sumout ;
wire \op_1~14 ;
wire \op_1~17_sumout ;
wire \op_1~18 ;
wire \op_1~21_sumout ;
wire \op_1~22 ;
wire \op_1~25_sumout ;
wire \op_1~26 ;
wire \op_1~29_sumout ;
wire \op_1~30 ;
wire \op_1~33_sumout ;
wire \op_1~34 ;
wire \op_1~37_sumout ;
wire \op_1~38 ;
wire \op_1~41_sumout ;
wire \op_1~42 ;
wire \op_1~45_sumout ;
wire \op_1~46 ;
wire \op_1~49_sumout ;
wire \op_1~50 ;
wire \op_1~53_sumout ;
wire \op_1~54 ;
wire \op_1~57_sumout ;
wire \op_1~58 ;
wire \op_1~61_sumout ;
wire \op_1~62 ;
wire \op_1~65_sumout ;
wire \op_1~66 ;
wire \op_1~69_sumout ;


dffeas \pipeline_dffe[0] (
	.clk(clock),
	.d(\op_1~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_0),
	.prn(vcc));
defparam \pipeline_dffe[0] .is_wysiwyg = "true";
defparam \pipeline_dffe[0] .power_up = "low";

dffeas \pipeline_dffe[1] (
	.clk(clock),
	.d(\op_1~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_1),
	.prn(vcc));
defparam \pipeline_dffe[1] .is_wysiwyg = "true";
defparam \pipeline_dffe[1] .power_up = "low";

dffeas \pipeline_dffe[2] (
	.clk(clock),
	.d(\op_1~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \pipeline_dffe[2] .is_wysiwyg = "true";
defparam \pipeline_dffe[2] .power_up = "low";

dffeas \pipeline_dffe[3] (
	.clk(clock),
	.d(\op_1~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \pipeline_dffe[3] .is_wysiwyg = "true";
defparam \pipeline_dffe[3] .power_up = "low";

dffeas \pipeline_dffe[4] (
	.clk(clock),
	.d(\op_1~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \pipeline_dffe[4] .is_wysiwyg = "true";
defparam \pipeline_dffe[4] .power_up = "low";

dffeas \pipeline_dffe[5] (
	.clk(clock),
	.d(\op_1~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \pipeline_dffe[5] .is_wysiwyg = "true";
defparam \pipeline_dffe[5] .power_up = "low";

dffeas \pipeline_dffe[6] (
	.clk(clock),
	.d(\op_1~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \pipeline_dffe[6] .is_wysiwyg = "true";
defparam \pipeline_dffe[6] .power_up = "low";

dffeas \pipeline_dffe[7] (
	.clk(clock),
	.d(\op_1~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \pipeline_dffe[7] .is_wysiwyg = "true";
defparam \pipeline_dffe[7] .power_up = "low";

dffeas \pipeline_dffe[8] (
	.clk(clock),
	.d(\op_1~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \pipeline_dffe[8] .is_wysiwyg = "true";
defparam \pipeline_dffe[8] .power_up = "low";

dffeas \pipeline_dffe[9] (
	.clk(clock),
	.d(\op_1~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \pipeline_dffe[9] .is_wysiwyg = "true";
defparam \pipeline_dffe[9] .power_up = "low";

dffeas \pipeline_dffe[10] (
	.clk(clock),
	.d(\op_1~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \pipeline_dffe[10] .is_wysiwyg = "true";
defparam \pipeline_dffe[10] .power_up = "low";

dffeas \pipeline_dffe[11] (
	.clk(clock),
	.d(\op_1~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \pipeline_dffe[11] .is_wysiwyg = "true";
defparam \pipeline_dffe[11] .power_up = "low";

dffeas \pipeline_dffe[12] (
	.clk(clock),
	.d(\op_1~49_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_12),
	.prn(vcc));
defparam \pipeline_dffe[12] .is_wysiwyg = "true";
defparam \pipeline_dffe[12] .power_up = "low";

dffeas \pipeline_dffe[13] (
	.clk(clock),
	.d(\op_1~53_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_13),
	.prn(vcc));
defparam \pipeline_dffe[13] .is_wysiwyg = "true";
defparam \pipeline_dffe[13] .power_up = "low";

dffeas \pipeline_dffe[14] (
	.clk(clock),
	.d(\op_1~57_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_14),
	.prn(vcc));
defparam \pipeline_dffe[14] .is_wysiwyg = "true";
defparam \pipeline_dffe[14] .power_up = "low";

dffeas \pipeline_dffe[15] (
	.clk(clock),
	.d(\op_1~61_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_15),
	.prn(vcc));
defparam \pipeline_dffe[15] .is_wysiwyg = "true";
defparam \pipeline_dffe[15] .power_up = "low";

dffeas \pipeline_dffe[16] (
	.clk(clock),
	.d(\op_1~65_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_16),
	.prn(vcc));
defparam \pipeline_dffe[16] .is_wysiwyg = "true";
defparam \pipeline_dffe[16] .power_up = "low";

dffeas \pipeline_dffe[17] (
	.clk(clock),
	.d(\op_1~69_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_17),
	.prn(vcc));
defparam \pipeline_dffe[17] .is_wysiwyg = "true";
defparam \pipeline_dffe[17] .power_up = "low";

arriav_lcell_comb \op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~1_sumout ),
	.cout(\op_1~2 ),
	.shareout());
defparam \op_1~1 .extended_lut = "off";
defparam \op_1~1 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~1 .shared_arith = "off";

arriav_lcell_comb \op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\op_1~2 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~5_sumout ),
	.cout(\op_1~6 ),
	.shareout());
defparam \op_1~5 .extended_lut = "off";
defparam \op_1~5 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~5 .shared_arith = "off";

arriav_lcell_comb \op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~9_sumout ),
	.cout(\op_1~10 ),
	.shareout());
defparam \op_1~9 .extended_lut = "off";
defparam \op_1~9 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~9 .shared_arith = "off";

arriav_lcell_comb \op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~13_sumout ),
	.cout(\op_1~14 ),
	.shareout());
defparam \op_1~13 .extended_lut = "off";
defparam \op_1~13 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~13 .shared_arith = "off";

arriav_lcell_comb \op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~17_sumout ),
	.cout(\op_1~18 ),
	.shareout());
defparam \op_1~17 .extended_lut = "off";
defparam \op_1~17 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~17 .shared_arith = "off";

arriav_lcell_comb \op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~21_sumout ),
	.cout(\op_1~22 ),
	.shareout());
defparam \op_1~21 .extended_lut = "off";
defparam \op_1~21 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~21 .shared_arith = "off";

arriav_lcell_comb \op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~25_sumout ),
	.cout(\op_1~26 ),
	.shareout());
defparam \op_1~25 .extended_lut = "off";
defparam \op_1~25 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~25 .shared_arith = "off";

arriav_lcell_comb \op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~29_sumout ),
	.cout(\op_1~30 ),
	.shareout());
defparam \op_1~29 .extended_lut = "off";
defparam \op_1~29 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~29 .shared_arith = "off";

arriav_lcell_comb \op_1~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\op_1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~33_sumout ),
	.cout(\op_1~34 ),
	.shareout());
defparam \op_1~33 .extended_lut = "off";
defparam \op_1~33 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~33 .shared_arith = "off";

arriav_lcell_comb \op_1~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\op_1~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~37_sumout ),
	.cout(\op_1~38 ),
	.shareout());
defparam \op_1~37 .extended_lut = "off";
defparam \op_1~37 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~37 .shared_arith = "off";

arriav_lcell_comb \op_1~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\op_1~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~41_sumout ),
	.cout(\op_1~42 ),
	.shareout());
defparam \op_1~41 .extended_lut = "off";
defparam \op_1~41 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~41 .shared_arith = "off";

arriav_lcell_comb \op_1~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\op_1~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~45_sumout ),
	.cout(\op_1~46 ),
	.shareout());
defparam \op_1~45 .extended_lut = "off";
defparam \op_1~45 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~45 .shared_arith = "off";

arriav_lcell_comb \op_1~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\op_1~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~49_sumout ),
	.cout(\op_1~50 ),
	.shareout());
defparam \op_1~49 .extended_lut = "off";
defparam \op_1~49 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~49 .shared_arith = "off";

arriav_lcell_comb \op_1~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\op_1~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~53_sumout ),
	.cout(\op_1~54 ),
	.shareout());
defparam \op_1~53 .extended_lut = "off";
defparam \op_1~53 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~53 .shared_arith = "off";

arriav_lcell_comb \op_1~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\op_1~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~57_sumout ),
	.cout(\op_1~58 ),
	.shareout());
defparam \op_1~57 .extended_lut = "off";
defparam \op_1~57 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~57 .shared_arith = "off";

arriav_lcell_comb \op_1~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\op_1~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~61_sumout ),
	.cout(\op_1~62 ),
	.shareout());
defparam \op_1~61 .extended_lut = "off";
defparam \op_1~61 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~61 .shared_arith = "off";

arriav_lcell_comb \op_1~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_16),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\op_1~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~65_sumout ),
	.cout(\op_1~66 ),
	.shareout());
defparam \op_1~65 .extended_lut = "off";
defparam \op_1~65 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~65 .shared_arith = "off";

arriav_lcell_comb \op_1~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_17),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\op_1~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~69_sumout ),
	.cout(),
	.shareout());
defparam \op_1~69 .extended_lut = "off";
defparam \op_1~69 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~69 .shared_arith = "off";

endmodule

module nco_test_lpm_add_sub_17 (
	a_0,
	xordvalue_11,
	a_10,
	pipeline_dffe_17,
	pipeline_dffe_16,
	pipeline_dffe_15,
	pipeline_dffe_14,
	pipeline_dffe_13,
	pipeline_dffe_12,
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_7,
	pipeline_dffe_6,
	pipeline_dffe_5,
	pipeline_dffe_4,
	pipeline_dffe_3,
	pipeline_dffe_2,
	pipeline_dffe_1,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_0;
input 	xordvalue_11;
input 	a_10;
output 	pipeline_dffe_17;
output 	pipeline_dffe_16;
output 	pipeline_dffe_15;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_7;
output 	pipeline_dffe_6;
output 	pipeline_dffe_5;
output 	pipeline_dffe_4;
output 	pipeline_dffe_3;
output 	pipeline_dffe_2;
output 	pipeline_dffe_1;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_add_sub_0qg_15 auto_generated(
	.a_0(a_0),
	.xordvalue_11(xordvalue_11),
	.a_10(a_10),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_1(pipeline_dffe_1),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module nco_test_add_sub_0qg_15 (
	a_0,
	xordvalue_11,
	a_10,
	pipeline_dffe_17,
	pipeline_dffe_16,
	pipeline_dffe_15,
	pipeline_dffe_14,
	pipeline_dffe_13,
	pipeline_dffe_12,
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_7,
	pipeline_dffe_6,
	pipeline_dffe_5,
	pipeline_dffe_4,
	pipeline_dffe_3,
	pipeline_dffe_2,
	pipeline_dffe_1,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_0;
input 	xordvalue_11;
input 	a_10;
output 	pipeline_dffe_17;
output 	pipeline_dffe_16;
output 	pipeline_dffe_15;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_7;
output 	pipeline_dffe_6;
output 	pipeline_dffe_5;
output 	pipeline_dffe_4;
output 	pipeline_dffe_3;
output 	pipeline_dffe_2;
output 	pipeline_dffe_1;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \op_1~0_combout ;
wire \op_1~1_combout ;
wire \op_1~2_combout ;
wire \op_1~3_combout ;
wire \op_1~4_combout ;
wire \op_1~5_combout ;
wire \op_1~6_combout ;
wire \op_1~7_combout ;
wire \op_1~8_combout ;


dffeas \pipeline_dffe[17] (
	.clk(clock),
	.d(\op_1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_17),
	.prn(vcc));
defparam \pipeline_dffe[17] .is_wysiwyg = "true";
defparam \pipeline_dffe[17] .power_up = "low";

dffeas \pipeline_dffe[16] (
	.clk(clock),
	.d(\op_1~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_16),
	.prn(vcc));
defparam \pipeline_dffe[16] .is_wysiwyg = "true";
defparam \pipeline_dffe[16] .power_up = "low";

dffeas \pipeline_dffe[15] (
	.clk(clock),
	.d(\op_1~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_15),
	.prn(vcc));
defparam \pipeline_dffe[15] .is_wysiwyg = "true";
defparam \pipeline_dffe[15] .power_up = "low";

dffeas \pipeline_dffe[14] (
	.clk(clock),
	.d(\op_1~3_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_14),
	.prn(vcc));
defparam \pipeline_dffe[14] .is_wysiwyg = "true";
defparam \pipeline_dffe[14] .power_up = "low";

dffeas \pipeline_dffe[13] (
	.clk(clock),
	.d(\op_1~4_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_13),
	.prn(vcc));
defparam \pipeline_dffe[13] .is_wysiwyg = "true";
defparam \pipeline_dffe[13] .power_up = "low";

dffeas \pipeline_dffe[12] (
	.clk(clock),
	.d(\op_1~5_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_12),
	.prn(vcc));
defparam \pipeline_dffe[12] .is_wysiwyg = "true";
defparam \pipeline_dffe[12] .power_up = "low";

dffeas \pipeline_dffe[11] (
	.clk(clock),
	.d(\op_1~6_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \pipeline_dffe[11] .is_wysiwyg = "true";
defparam \pipeline_dffe[11] .power_up = "low";

dffeas \pipeline_dffe[10] (
	.clk(clock),
	.d(\op_1~4_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \pipeline_dffe[10] .is_wysiwyg = "true";
defparam \pipeline_dffe[10] .power_up = "low";

dffeas \pipeline_dffe[9] (
	.clk(clock),
	.d(\op_1~5_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \pipeline_dffe[9] .is_wysiwyg = "true";
defparam \pipeline_dffe[9] .power_up = "low";

dffeas \pipeline_dffe[8] (
	.clk(clock),
	.d(\op_1~6_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \pipeline_dffe[8] .is_wysiwyg = "true";
defparam \pipeline_dffe[8] .power_up = "low";

dffeas \pipeline_dffe[7] (
	.clk(clock),
	.d(\op_1~4_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \pipeline_dffe[7] .is_wysiwyg = "true";
defparam \pipeline_dffe[7] .power_up = "low";

dffeas \pipeline_dffe[6] (
	.clk(clock),
	.d(\op_1~5_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \pipeline_dffe[6] .is_wysiwyg = "true";
defparam \pipeline_dffe[6] .power_up = "low";

dffeas \pipeline_dffe[5] (
	.clk(clock),
	.d(\op_1~7_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \pipeline_dffe[5] .is_wysiwyg = "true";
defparam \pipeline_dffe[5] .power_up = "low";

dffeas \pipeline_dffe[4] (
	.clk(clock),
	.d(\op_1~2_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \pipeline_dffe[4] .is_wysiwyg = "true";
defparam \pipeline_dffe[4] .power_up = "low";

dffeas \pipeline_dffe[3] (
	.clk(clock),
	.d(\op_1~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \pipeline_dffe[3] .is_wysiwyg = "true";
defparam \pipeline_dffe[3] .power_up = "low";

dffeas \pipeline_dffe[2] (
	.clk(clock),
	.d(\op_1~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \pipeline_dffe[2] .is_wysiwyg = "true";
defparam \pipeline_dffe[2] .power_up = "low";

dffeas \pipeline_dffe[1] (
	.clk(clock),
	.d(\op_1~8_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_1),
	.prn(vcc));
defparam \pipeline_dffe[1] .is_wysiwyg = "true";
defparam \pipeline_dffe[1] .power_up = "low";

arriav_lcell_comb \op_1~0 (
	.dataa(!a_0),
	.datab(!xordvalue_11),
	.datac(!a_10),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\op_1~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \op_1~0 .extended_lut = "off";
defparam \op_1~0 .lut_mask = 64'hFDFDFDFDFDFDFDFD;
defparam \op_1~0 .shared_arith = "off";

arriav_lcell_comb \op_1~1 (
	.dataa(!a_0),
	.datab(!xordvalue_11),
	.datac(!a_10),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\op_1~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \op_1~1 .extended_lut = "off";
defparam \op_1~1 .lut_mask = 64'h9696969696969696;
defparam \op_1~1 .shared_arith = "off";

arriav_lcell_comb \op_1~2 (
	.dataa(!a_0),
	.datab(!xordvalue_11),
	.datac(!a_10),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\op_1~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \op_1~2 .extended_lut = "off";
defparam \op_1~2 .lut_mask = 64'h6F6F6F6F6F6F6F6F;
defparam \op_1~2 .shared_arith = "off";

arriav_lcell_comb \op_1~3 (
	.dataa(!a_0),
	.datab(!xordvalue_11),
	.datac(!a_10),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\op_1~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \op_1~3 .extended_lut = "off";
defparam \op_1~3 .lut_mask = 64'h9696969696969696;
defparam \op_1~3 .shared_arith = "off";

arriav_lcell_comb \op_1~4 (
	.dataa(!a_0),
	.datab(!xordvalue_11),
	.datac(!a_10),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\op_1~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \op_1~4 .extended_lut = "off";
defparam \op_1~4 .lut_mask = 64'h9696969696969696;
defparam \op_1~4 .shared_arith = "off";

arriav_lcell_comb \op_1~5 (
	.dataa(!a_0),
	.datab(!xordvalue_11),
	.datac(!a_10),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\op_1~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \op_1~5 .extended_lut = "off";
defparam \op_1~5 .lut_mask = 64'hBFBFBFBFBFBFBFBF;
defparam \op_1~5 .shared_arith = "off";

arriav_lcell_comb \op_1~6 (
	.dataa(!a_0),
	.datab(!xordvalue_11),
	.datac(!a_10),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\op_1~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \op_1~6 .extended_lut = "off";
defparam \op_1~6 .lut_mask = 64'h9696969696969696;
defparam \op_1~6 .shared_arith = "off";

arriav_lcell_comb \op_1~7 (
	.dataa(!a_0),
	.datab(!xordvalue_11),
	.datac(!a_10),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\op_1~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \op_1~7 .extended_lut = "off";
defparam \op_1~7 .lut_mask = 64'h9696969696969696;
defparam \op_1~7 .shared_arith = "off";

arriav_lcell_comb \op_1~8 (
	.dataa(!a_0),
	.datab(!xordvalue_11),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\op_1~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \op_1~8 .extended_lut = "off";
defparam \op_1~8 .lut_mask = 64'h6666666666666666;
defparam \op_1~8 .shared_arith = "off";

endmodule

module nco_test_cordic_axor_1p_lpm_16 (
	sin_o_0,
	pipeline_dffe_17,
	pipeline_dffe_16,
	dffe16,
	pipeline_dffe_15,
	pipeline_dffe_171,
	dffe18,
	pipeline_dffe_14,
	pipeline_dffe_161,
	pipeline_dffe_13,
	dffe17,
	pipeline_dffe_151,
	pipeline_dffe_12,
	dffe161,
	pipeline_dffe_141,
	pipeline_dffe_11,
	dffe15,
	pipeline_dffe_131,
	pipeline_dffe_10,
	dffe14,
	pipeline_dffe_121,
	pipeline_dffe_9,
	dffe13,
	pipeline_dffe_111,
	pipeline_dffe_8,
	dffe12,
	pipeline_dffe_101,
	pipeline_dffe_7,
	dffe11,
	pipeline_dffe_91,
	pipeline_dffe_6,
	dffe10,
	pipeline_dffe_81,
	pipeline_dffe_5,
	dffe9,
	pipeline_dffe_71,
	pipeline_dffe_4,
	dffe8,
	pipeline_dffe_3,
	pipeline_dffe_61,
	pipeline_dffe_0,
	dffe7,
	pipeline_dffe_51,
	pipeline_dffe_1,
	pipeline_dffe_2,
	dffe6,
	pipeline_dffe_41,
	dffe5,
	pipeline_dffe_31,
	dffe3,
	dffe4,
	pipeline_dffe_21,
	pipeline_dffe_18,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	sin_o_0;
output 	pipeline_dffe_17;
output 	pipeline_dffe_16;
input 	dffe16;
output 	pipeline_dffe_15;
input 	pipeline_dffe_171;
input 	dffe18;
output 	pipeline_dffe_14;
input 	pipeline_dffe_161;
output 	pipeline_dffe_13;
input 	dffe17;
input 	pipeline_dffe_151;
output 	pipeline_dffe_12;
input 	dffe161;
input 	pipeline_dffe_141;
output 	pipeline_dffe_11;
input 	dffe15;
input 	pipeline_dffe_131;
output 	pipeline_dffe_10;
input 	dffe14;
input 	pipeline_dffe_121;
output 	pipeline_dffe_9;
input 	dffe13;
input 	pipeline_dffe_111;
output 	pipeline_dffe_8;
input 	dffe12;
input 	pipeline_dffe_101;
output 	pipeline_dffe_7;
input 	dffe11;
input 	pipeline_dffe_91;
output 	pipeline_dffe_6;
input 	dffe10;
input 	pipeline_dffe_81;
output 	pipeline_dffe_5;
input 	dffe9;
input 	pipeline_dffe_71;
output 	pipeline_dffe_4;
input 	dffe8;
output 	pipeline_dffe_3;
input 	pipeline_dffe_61;
output 	pipeline_dffe_0;
input 	dffe7;
input 	pipeline_dffe_51;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
input 	dffe6;
input 	pipeline_dffe_41;
input 	dffe5;
input 	pipeline_dffe_31;
input 	dffe3;
input 	dffe4;
input 	pipeline_dffe_21;
input 	pipeline_dffe_18;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[17]~q ;
wire \xordvalue[15]~q ;
wire \a[16]~q ;
wire \a[15]~q ;
wire \a[14]~q ;
wire \xordvalue[14]~q ;
wire \a[13]~q ;
wire \xordvalue[13]~q ;
wire \a[12]~q ;
wire \xordvalue[12]~q ;
wire \a[11]~q ;
wire \xordvalue[11]~q ;
wire \a[10]~q ;
wire \xordvalue[10]~q ;
wire \a[9]~q ;
wire \xordvalue[9]~q ;
wire \a[8]~q ;
wire \xordvalue[8]~q ;
wire \a[7]~q ;
wire \xordvalue[7]~q ;
wire \a[6]~q ;
wire \xordvalue[6]~q ;
wire \a[5]~q ;
wire \xordvalue[5]~q ;
wire \a[4]~q ;
wire \xordvalue[4]~q ;
wire \a[3]~q ;
wire \xordvalue[3]~q ;
wire \a[0]~q ;
wire \xordvalue[0]~q ;
wire \a[2]~q ;
wire \xordvalue[2]~q ;
wire \a[1]~q ;
wire \xordvalue[1]~q ;
wire \xordvalue~0_combout ;
wire \xordvalue~1_combout ;
wire \xordvalue~2_combout ;
wire \xordvalue~3_combout ;
wire \xordvalue~4_combout ;
wire \xordvalue~5_combout ;
wire \xordvalue~6_combout ;
wire \xordvalue~7_combout ;
wire \xordvalue~8_combout ;
wire \xordvalue~9_combout ;
wire \xordvalue~10_combout ;
wire \xordvalue~11_combout ;
wire \xordvalue~12_combout ;
wire \xordvalue~13_combout ;
wire \xordvalue~14_combout ;
wire \xordvalue~15_combout ;


nco_test_lpm_add_sub_18 u0(
	.a_17(\a[17]~q ),
	.xordvalue_15(\xordvalue[15]~q ),
	.a_16(\a[16]~q ),
	.a_15(\a[15]~q ),
	.a_14(\a[14]~q ),
	.xordvalue_14(\xordvalue[14]~q ),
	.a_13(\a[13]~q ),
	.xordvalue_13(\xordvalue[13]~q ),
	.a_12(\a[12]~q ),
	.xordvalue_12(\xordvalue[12]~q ),
	.a_11(\a[11]~q ),
	.xordvalue_11(\xordvalue[11]~q ),
	.a_10(\a[10]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.a_9(\a[9]~q ),
	.xordvalue_9(\xordvalue[9]~q ),
	.a_8(\a[8]~q ),
	.xordvalue_8(\xordvalue[8]~q ),
	.a_7(\a[7]~q ),
	.xordvalue_7(\xordvalue[7]~q ),
	.a_6(\a[6]~q ),
	.xordvalue_6(\xordvalue[6]~q ),
	.a_5(\a[5]~q ),
	.xordvalue_5(\xordvalue[5]~q ),
	.a_4(\a[4]~q ),
	.xordvalue_4(\xordvalue[4]~q ),
	.a_3(\a[3]~q ),
	.xordvalue_3(\xordvalue[3]~q ),
	.a_0(\a[0]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_2(\a[2]~q ),
	.xordvalue_2(\xordvalue[2]~q ),
	.a_1(\a[1]~q ),
	.xordvalue_1(\xordvalue[1]~q ),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[17] (
	.clk(clk),
	.d(pipeline_dffe_171),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[17]~q ),
	.prn(vcc));
defparam \a[17] .is_wysiwyg = "true";
defparam \a[17] .power_up = "low";

dffeas \xordvalue[15] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[15]~q ),
	.prn(vcc));
defparam \xordvalue[15] .is_wysiwyg = "true";
defparam \xordvalue[15] .power_up = "low";

dffeas \a[16] (
	.clk(clk),
	.d(pipeline_dffe_161),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[16]~q ),
	.prn(vcc));
defparam \a[16] .is_wysiwyg = "true";
defparam \a[16] .power_up = "low";

dffeas \a[15] (
	.clk(clk),
	.d(pipeline_dffe_151),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

dffeas \a[14] (
	.clk(clk),
	.d(pipeline_dffe_141),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

dffeas \xordvalue[14] (
	.clk(clk),
	.d(\xordvalue~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[14]~q ),
	.prn(vcc));
defparam \xordvalue[14] .is_wysiwyg = "true";
defparam \xordvalue[14] .power_up = "low";

dffeas \a[13] (
	.clk(clk),
	.d(pipeline_dffe_131),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

dffeas \xordvalue[13] (
	.clk(clk),
	.d(\xordvalue~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[13]~q ),
	.prn(vcc));
defparam \xordvalue[13] .is_wysiwyg = "true";
defparam \xordvalue[13] .power_up = "low";

dffeas \a[12] (
	.clk(clk),
	.d(pipeline_dffe_121),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

dffeas \xordvalue[12] (
	.clk(clk),
	.d(\xordvalue~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[12]~q ),
	.prn(vcc));
defparam \xordvalue[12] .is_wysiwyg = "true";
defparam \xordvalue[12] .power_up = "low";

dffeas \a[11] (
	.clk(clk),
	.d(pipeline_dffe_111),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \xordvalue[11] (
	.clk(clk),
	.d(\xordvalue~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[11]~q ),
	.prn(vcc));
defparam \xordvalue[11] .is_wysiwyg = "true";
defparam \xordvalue[11] .power_up = "low";

dffeas \a[10] (
	.clk(clk),
	.d(pipeline_dffe_101),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(\xordvalue~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

dffeas \a[9] (
	.clk(clk),
	.d(pipeline_dffe_91),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \xordvalue[9] (
	.clk(clk),
	.d(\xordvalue~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[9]~q ),
	.prn(vcc));
defparam \xordvalue[9] .is_wysiwyg = "true";
defparam \xordvalue[9] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(pipeline_dffe_81),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \xordvalue[8] (
	.clk(clk),
	.d(\xordvalue~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[8]~q ),
	.prn(vcc));
defparam \xordvalue[8] .is_wysiwyg = "true";
defparam \xordvalue[8] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(pipeline_dffe_71),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \xordvalue[7] (
	.clk(clk),
	.d(\xordvalue~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[7]~q ),
	.prn(vcc));
defparam \xordvalue[7] .is_wysiwyg = "true";
defparam \xordvalue[7] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(pipeline_dffe_61),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \xordvalue[6] (
	.clk(clk),
	.d(\xordvalue~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[6]~q ),
	.prn(vcc));
defparam \xordvalue[6] .is_wysiwyg = "true";
defparam \xordvalue[6] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(pipeline_dffe_51),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \xordvalue[5] (
	.clk(clk),
	.d(\xordvalue~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[5]~q ),
	.prn(vcc));
defparam \xordvalue[5] .is_wysiwyg = "true";
defparam \xordvalue[5] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(pipeline_dffe_41),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \xordvalue[4] (
	.clk(clk),
	.d(\xordvalue~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[4]~q ),
	.prn(vcc));
defparam \xordvalue[4] .is_wysiwyg = "true";
defparam \xordvalue[4] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(pipeline_dffe_31),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \xordvalue[3] (
	.clk(clk),
	.d(\xordvalue~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[3]~q ),
	.prn(vcc));
defparam \xordvalue[3] .is_wysiwyg = "true";
defparam \xordvalue[3] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(dffe16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(pipeline_dffe_21),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \xordvalue[2] (
	.clk(clk),
	.d(\xordvalue~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[2]~q ),
	.prn(vcc));
defparam \xordvalue[2] .is_wysiwyg = "true";
defparam \xordvalue[2] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(pipeline_dffe_18),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \xordvalue[1] (
	.clk(clk),
	.d(\xordvalue~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[1]~q ),
	.prn(vcc));
defparam \xordvalue[1] .is_wysiwyg = "true";
defparam \xordvalue[1] .power_up = "low";

arriav_lcell_comb \xordvalue~0 (
	.dataa(!dffe18),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

arriav_lcell_comb \xordvalue~1 (
	.dataa(!dffe17),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~1 .extended_lut = "off";
defparam \xordvalue~1 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~1 .shared_arith = "off";

arriav_lcell_comb \xordvalue~2 (
	.dataa(!dffe161),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~2 .extended_lut = "off";
defparam \xordvalue~2 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~2 .shared_arith = "off";

arriav_lcell_comb \xordvalue~3 (
	.dataa(!dffe15),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~3 .extended_lut = "off";
defparam \xordvalue~3 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~3 .shared_arith = "off";

arriav_lcell_comb \xordvalue~4 (
	.dataa(!dffe14),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~4 .extended_lut = "off";
defparam \xordvalue~4 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~4 .shared_arith = "off";

arriav_lcell_comb \xordvalue~5 (
	.dataa(!dffe13),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~5 .extended_lut = "off";
defparam \xordvalue~5 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~5 .shared_arith = "off";

arriav_lcell_comb \xordvalue~6 (
	.dataa(!dffe12),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~6 .extended_lut = "off";
defparam \xordvalue~6 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~6 .shared_arith = "off";

arriav_lcell_comb \xordvalue~7 (
	.dataa(!dffe11),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~7 .extended_lut = "off";
defparam \xordvalue~7 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~7 .shared_arith = "off";

arriav_lcell_comb \xordvalue~8 (
	.dataa(!dffe10),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~8 .extended_lut = "off";
defparam \xordvalue~8 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~8 .shared_arith = "off";

arriav_lcell_comb \xordvalue~9 (
	.dataa(!dffe9),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~9 .extended_lut = "off";
defparam \xordvalue~9 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~9 .shared_arith = "off";

arriav_lcell_comb \xordvalue~10 (
	.dataa(!dffe8),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~10 .extended_lut = "off";
defparam \xordvalue~10 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~10 .shared_arith = "off";

arriav_lcell_comb \xordvalue~11 (
	.dataa(!dffe7),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~11 .extended_lut = "off";
defparam \xordvalue~11 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~11 .shared_arith = "off";

arriav_lcell_comb \xordvalue~12 (
	.dataa(!dffe6),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~12 .extended_lut = "off";
defparam \xordvalue~12 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~12 .shared_arith = "off";

arriav_lcell_comb \xordvalue~13 (
	.dataa(!dffe3),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~13 .extended_lut = "off";
defparam \xordvalue~13 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~13 .shared_arith = "off";

arriav_lcell_comb \xordvalue~14 (
	.dataa(!dffe5),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~14 .extended_lut = "off";
defparam \xordvalue~14 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~14 .shared_arith = "off";

arriav_lcell_comb \xordvalue~15 (
	.dataa(!dffe4),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~15 .extended_lut = "off";
defparam \xordvalue~15 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~15 .shared_arith = "off";

endmodule

module nco_test_lpm_add_sub_18 (
	a_17,
	xordvalue_15,
	a_16,
	a_15,
	a_14,
	xordvalue_14,
	a_13,
	xordvalue_13,
	a_12,
	xordvalue_12,
	a_11,
	xordvalue_11,
	a_10,
	xordvalue_10,
	a_9,
	xordvalue_9,
	a_8,
	xordvalue_8,
	a_7,
	xordvalue_7,
	a_6,
	xordvalue_6,
	a_5,
	xordvalue_5,
	a_4,
	xordvalue_4,
	a_3,
	xordvalue_3,
	a_0,
	xordvalue_0,
	a_2,
	xordvalue_2,
	a_1,
	xordvalue_1,
	pipeline_dffe_17,
	pipeline_dffe_16,
	pipeline_dffe_15,
	pipeline_dffe_14,
	pipeline_dffe_13,
	pipeline_dffe_12,
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_7,
	pipeline_dffe_6,
	pipeline_dffe_5,
	pipeline_dffe_4,
	pipeline_dffe_3,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_15;
input 	a_16;
input 	a_15;
input 	a_14;
input 	xordvalue_14;
input 	a_13;
input 	xordvalue_13;
input 	a_12;
input 	xordvalue_12;
input 	a_11;
input 	xordvalue_11;
input 	a_10;
input 	xordvalue_10;
input 	a_9;
input 	xordvalue_9;
input 	a_8;
input 	xordvalue_8;
input 	a_7;
input 	xordvalue_7;
input 	a_6;
input 	xordvalue_6;
input 	a_5;
input 	xordvalue_5;
input 	a_4;
input 	xordvalue_4;
input 	a_3;
input 	xordvalue_3;
input 	a_0;
input 	xordvalue_0;
input 	a_2;
input 	xordvalue_2;
input 	a_1;
input 	xordvalue_1;
output 	pipeline_dffe_17;
output 	pipeline_dffe_16;
output 	pipeline_dffe_15;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_7;
output 	pipeline_dffe_6;
output 	pipeline_dffe_5;
output 	pipeline_dffe_4;
output 	pipeline_dffe_3;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_add_sub_0qg_16 auto_generated(
	.a_17(a_17),
	.xordvalue_15(xordvalue_15),
	.a_16(a_16),
	.a_15(a_15),
	.a_14(a_14),
	.xordvalue_14(xordvalue_14),
	.a_13(a_13),
	.xordvalue_13(xordvalue_13),
	.a_12(a_12),
	.xordvalue_12(xordvalue_12),
	.a_11(a_11),
	.xordvalue_11(xordvalue_11),
	.a_10(a_10),
	.xordvalue_10(xordvalue_10),
	.a_9(a_9),
	.xordvalue_9(xordvalue_9),
	.a_8(a_8),
	.xordvalue_8(xordvalue_8),
	.a_7(a_7),
	.xordvalue_7(xordvalue_7),
	.a_6(a_6),
	.xordvalue_6(xordvalue_6),
	.a_5(a_5),
	.xordvalue_5(xordvalue_5),
	.a_4(a_4),
	.xordvalue_4(xordvalue_4),
	.a_3(a_3),
	.xordvalue_3(xordvalue_3),
	.a_0(a_0),
	.xordvalue_0(xordvalue_0),
	.a_2(a_2),
	.xordvalue_2(xordvalue_2),
	.a_1(a_1),
	.xordvalue_1(xordvalue_1),
	.pipeline_dffe_17(pipeline_dffe_17),
	.pipeline_dffe_16(pipeline_dffe_16),
	.pipeline_dffe_15(pipeline_dffe_15),
	.pipeline_dffe_14(pipeline_dffe_14),
	.pipeline_dffe_13(pipeline_dffe_13),
	.pipeline_dffe_12(pipeline_dffe_12),
	.pipeline_dffe_11(pipeline_dffe_11),
	.pipeline_dffe_10(pipeline_dffe_10),
	.pipeline_dffe_9(pipeline_dffe_9),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_2(pipeline_dffe_2),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module nco_test_add_sub_0qg_16 (
	a_17,
	xordvalue_15,
	a_16,
	a_15,
	a_14,
	xordvalue_14,
	a_13,
	xordvalue_13,
	a_12,
	xordvalue_12,
	a_11,
	xordvalue_11,
	a_10,
	xordvalue_10,
	a_9,
	xordvalue_9,
	a_8,
	xordvalue_8,
	a_7,
	xordvalue_7,
	a_6,
	xordvalue_6,
	a_5,
	xordvalue_5,
	a_4,
	xordvalue_4,
	a_3,
	xordvalue_3,
	a_0,
	xordvalue_0,
	a_2,
	xordvalue_2,
	a_1,
	xordvalue_1,
	pipeline_dffe_17,
	pipeline_dffe_16,
	pipeline_dffe_15,
	pipeline_dffe_14,
	pipeline_dffe_13,
	pipeline_dffe_12,
	pipeline_dffe_11,
	pipeline_dffe_10,
	pipeline_dffe_9,
	pipeline_dffe_8,
	pipeline_dffe_7,
	pipeline_dffe_6,
	pipeline_dffe_5,
	pipeline_dffe_4,
	pipeline_dffe_3,
	pipeline_dffe_0,
	pipeline_dffe_1,
	pipeline_dffe_2,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_15;
input 	a_16;
input 	a_15;
input 	a_14;
input 	xordvalue_14;
input 	a_13;
input 	xordvalue_13;
input 	a_12;
input 	xordvalue_12;
input 	a_11;
input 	xordvalue_11;
input 	a_10;
input 	xordvalue_10;
input 	a_9;
input 	xordvalue_9;
input 	a_8;
input 	xordvalue_8;
input 	a_7;
input 	xordvalue_7;
input 	a_6;
input 	xordvalue_6;
input 	a_5;
input 	xordvalue_5;
input 	a_4;
input 	xordvalue_4;
input 	a_3;
input 	xordvalue_3;
input 	a_0;
input 	xordvalue_0;
input 	a_2;
input 	xordvalue_2;
input 	a_1;
input 	xordvalue_1;
output 	pipeline_dffe_17;
output 	pipeline_dffe_16;
output 	pipeline_dffe_15;
output 	pipeline_dffe_14;
output 	pipeline_dffe_13;
output 	pipeline_dffe_12;
output 	pipeline_dffe_11;
output 	pipeline_dffe_10;
output 	pipeline_dffe_9;
output 	pipeline_dffe_8;
output 	pipeline_dffe_7;
output 	pipeline_dffe_6;
output 	pipeline_dffe_5;
output 	pipeline_dffe_4;
output 	pipeline_dffe_3;
output 	pipeline_dffe_0;
output 	pipeline_dffe_1;
output 	pipeline_dffe_2;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \op_1~62 ;
wire \op_1~70 ;
wire \op_1~66 ;
wire \op_1~58 ;
wire \op_1~54 ;
wire \op_1~50 ;
wire \op_1~46 ;
wire \op_1~42 ;
wire \op_1~38 ;
wire \op_1~34 ;
wire \op_1~30 ;
wire \op_1~26 ;
wire \op_1~22 ;
wire \op_1~18 ;
wire \op_1~14 ;
wire \op_1~10 ;
wire \op_1~6 ;
wire \op_1~1_sumout ;
wire \op_1~5_sumout ;
wire \op_1~9_sumout ;
wire \op_1~13_sumout ;
wire \op_1~17_sumout ;
wire \op_1~21_sumout ;
wire \op_1~25_sumout ;
wire \op_1~29_sumout ;
wire \op_1~33_sumout ;
wire \op_1~37_sumout ;
wire \op_1~41_sumout ;
wire \op_1~45_sumout ;
wire \op_1~49_sumout ;
wire \op_1~53_sumout ;
wire \op_1~57_sumout ;
wire \op_1~61_sumout ;
wire \op_1~69_sumout ;
wire \op_1~65_sumout ;


dffeas \pipeline_dffe[17] (
	.clk(clock),
	.d(\op_1~1_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_17),
	.prn(vcc));
defparam \pipeline_dffe[17] .is_wysiwyg = "true";
defparam \pipeline_dffe[17] .power_up = "low";

dffeas \pipeline_dffe[16] (
	.clk(clock),
	.d(\op_1~5_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_16),
	.prn(vcc));
defparam \pipeline_dffe[16] .is_wysiwyg = "true";
defparam \pipeline_dffe[16] .power_up = "low";

dffeas \pipeline_dffe[15] (
	.clk(clock),
	.d(\op_1~9_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_15),
	.prn(vcc));
defparam \pipeline_dffe[15] .is_wysiwyg = "true";
defparam \pipeline_dffe[15] .power_up = "low";

dffeas \pipeline_dffe[14] (
	.clk(clock),
	.d(\op_1~13_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_14),
	.prn(vcc));
defparam \pipeline_dffe[14] .is_wysiwyg = "true";
defparam \pipeline_dffe[14] .power_up = "low";

dffeas \pipeline_dffe[13] (
	.clk(clock),
	.d(\op_1~17_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_13),
	.prn(vcc));
defparam \pipeline_dffe[13] .is_wysiwyg = "true";
defparam \pipeline_dffe[13] .power_up = "low";

dffeas \pipeline_dffe[12] (
	.clk(clock),
	.d(\op_1~21_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_12),
	.prn(vcc));
defparam \pipeline_dffe[12] .is_wysiwyg = "true";
defparam \pipeline_dffe[12] .power_up = "low";

dffeas \pipeline_dffe[11] (
	.clk(clock),
	.d(\op_1~25_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_11),
	.prn(vcc));
defparam \pipeline_dffe[11] .is_wysiwyg = "true";
defparam \pipeline_dffe[11] .power_up = "low";

dffeas \pipeline_dffe[10] (
	.clk(clock),
	.d(\op_1~29_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_10),
	.prn(vcc));
defparam \pipeline_dffe[10] .is_wysiwyg = "true";
defparam \pipeline_dffe[10] .power_up = "low";

dffeas \pipeline_dffe[9] (
	.clk(clock),
	.d(\op_1~33_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \pipeline_dffe[9] .is_wysiwyg = "true";
defparam \pipeline_dffe[9] .power_up = "low";

dffeas \pipeline_dffe[8] (
	.clk(clock),
	.d(\op_1~37_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \pipeline_dffe[8] .is_wysiwyg = "true";
defparam \pipeline_dffe[8] .power_up = "low";

dffeas \pipeline_dffe[7] (
	.clk(clock),
	.d(\op_1~41_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \pipeline_dffe[7] .is_wysiwyg = "true";
defparam \pipeline_dffe[7] .power_up = "low";

dffeas \pipeline_dffe[6] (
	.clk(clock),
	.d(\op_1~45_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \pipeline_dffe[6] .is_wysiwyg = "true";
defparam \pipeline_dffe[6] .power_up = "low";

dffeas \pipeline_dffe[5] (
	.clk(clock),
	.d(\op_1~49_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \pipeline_dffe[5] .is_wysiwyg = "true";
defparam \pipeline_dffe[5] .power_up = "low";

dffeas \pipeline_dffe[4] (
	.clk(clock),
	.d(\op_1~53_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \pipeline_dffe[4] .is_wysiwyg = "true";
defparam \pipeline_dffe[4] .power_up = "low";

dffeas \pipeline_dffe[3] (
	.clk(clock),
	.d(\op_1~57_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \pipeline_dffe[3] .is_wysiwyg = "true";
defparam \pipeline_dffe[3] .power_up = "low";

dffeas \pipeline_dffe[0] (
	.clk(clock),
	.d(\op_1~61_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_0),
	.prn(vcc));
defparam \pipeline_dffe[0] .is_wysiwyg = "true";
defparam \pipeline_dffe[0] .power_up = "low";

dffeas \pipeline_dffe[1] (
	.clk(clock),
	.d(\op_1~69_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_1),
	.prn(vcc));
defparam \pipeline_dffe[1] .is_wysiwyg = "true";
defparam \pipeline_dffe[1] .power_up = "low";

dffeas \pipeline_dffe[2] (
	.clk(clock),
	.d(\op_1~65_sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \pipeline_dffe[2] .is_wysiwyg = "true";
defparam \pipeline_dffe[2] .power_up = "low";

arriav_lcell_comb \op_1~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~61_sumout ),
	.cout(\op_1~62 ),
	.shareout());
defparam \op_1~61 .extended_lut = "off";
defparam \op_1~61 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~61 .shared_arith = "off";

arriav_lcell_comb \op_1~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_1),
	.datag(gnd),
	.cin(\op_1~62 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~69_sumout ),
	.cout(\op_1~70 ),
	.shareout());
defparam \op_1~69 .extended_lut = "off";
defparam \op_1~69 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~69 .shared_arith = "off";

arriav_lcell_comb \op_1~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_2),
	.datag(gnd),
	.cin(\op_1~70 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~65_sumout ),
	.cout(\op_1~66 ),
	.shareout());
defparam \op_1~65 .extended_lut = "off";
defparam \op_1~65 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~65 .shared_arith = "off";

arriav_lcell_comb \op_1~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_3),
	.datag(gnd),
	.cin(\op_1~66 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~57_sumout ),
	.cout(\op_1~58 ),
	.shareout());
defparam \op_1~57 .extended_lut = "off";
defparam \op_1~57 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~57 .shared_arith = "off";

arriav_lcell_comb \op_1~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_4),
	.datag(gnd),
	.cin(\op_1~58 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~53_sumout ),
	.cout(\op_1~54 ),
	.shareout());
defparam \op_1~53 .extended_lut = "off";
defparam \op_1~53 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~53 .shared_arith = "off";

arriav_lcell_comb \op_1~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_5),
	.datag(gnd),
	.cin(\op_1~54 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~49_sumout ),
	.cout(\op_1~50 ),
	.shareout());
defparam \op_1~49 .extended_lut = "off";
defparam \op_1~49 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~49 .shared_arith = "off";

arriav_lcell_comb \op_1~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_6),
	.datag(gnd),
	.cin(\op_1~50 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~45_sumout ),
	.cout(\op_1~46 ),
	.shareout());
defparam \op_1~45 .extended_lut = "off";
defparam \op_1~45 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~45 .shared_arith = "off";

arriav_lcell_comb \op_1~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_7),
	.datag(gnd),
	.cin(\op_1~46 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~41_sumout ),
	.cout(\op_1~42 ),
	.shareout());
defparam \op_1~41 .extended_lut = "off";
defparam \op_1~41 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~41 .shared_arith = "off";

arriav_lcell_comb \op_1~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_8),
	.datag(gnd),
	.cin(\op_1~42 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~37_sumout ),
	.cout(\op_1~38 ),
	.shareout());
defparam \op_1~37 .extended_lut = "off";
defparam \op_1~37 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~37 .shared_arith = "off";

arriav_lcell_comb \op_1~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_9),
	.datag(gnd),
	.cin(\op_1~38 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~33_sumout ),
	.cout(\op_1~34 ),
	.shareout());
defparam \op_1~33 .extended_lut = "off";
defparam \op_1~33 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~33 .shared_arith = "off";

arriav_lcell_comb \op_1~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\op_1~34 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~29_sumout ),
	.cout(\op_1~30 ),
	.shareout());
defparam \op_1~29 .extended_lut = "off";
defparam \op_1~29 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~29 .shared_arith = "off";

arriav_lcell_comb \op_1~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_11),
	.datag(gnd),
	.cin(\op_1~30 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~25_sumout ),
	.cout(\op_1~26 ),
	.shareout());
defparam \op_1~25 .extended_lut = "off";
defparam \op_1~25 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~25 .shared_arith = "off";

arriav_lcell_comb \op_1~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_12),
	.datag(gnd),
	.cin(\op_1~26 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~21_sumout ),
	.cout(\op_1~22 ),
	.shareout());
defparam \op_1~21 .extended_lut = "off";
defparam \op_1~21 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~21 .shared_arith = "off";

arriav_lcell_comb \op_1~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_13),
	.datag(gnd),
	.cin(\op_1~22 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~17_sumout ),
	.cout(\op_1~18 ),
	.shareout());
defparam \op_1~17 .extended_lut = "off";
defparam \op_1~17 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~17 .shared_arith = "off";

arriav_lcell_comb \op_1~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_14),
	.datag(gnd),
	.cin(\op_1~18 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~13_sumout ),
	.cout(\op_1~14 ),
	.shareout());
defparam \op_1~13 .extended_lut = "off";
defparam \op_1~13 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~13 .shared_arith = "off";

arriav_lcell_comb \op_1~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_15),
	.datag(gnd),
	.cin(\op_1~14 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~9_sumout ),
	.cout(\op_1~10 ),
	.shareout());
defparam \op_1~9 .extended_lut = "off";
defparam \op_1~9 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~9 .shared_arith = "off";

arriav_lcell_comb \op_1~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_16),
	.datae(gnd),
	.dataf(!xordvalue_15),
	.datag(gnd),
	.cin(\op_1~10 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~5_sumout ),
	.cout(\op_1~6 ),
	.shareout());
defparam \op_1~5 .extended_lut = "off";
defparam \op_1~5 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~5 .shared_arith = "off";

arriav_lcell_comb \op_1~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_17),
	.datae(gnd),
	.dataf(!xordvalue_15),
	.datag(gnd),
	.cin(\op_1~6 ),
	.sharein(gnd),
	.combout(),
	.sumout(\op_1~1_sumout ),
	.cout(),
	.shareout());
defparam \op_1~1 .extended_lut = "off";
defparam \op_1~1 .lut_mask = 64'h0000FF00000000FF;
defparam \op_1~1 .shared_arith = "off";

endmodule

module nco_test_cordic_sxor_1p_lpm (
	sin_o_0,
	dffe18,
	dffe17,
	dffe16,
	dffe161,
	dffe181,
	pipeline_dffe_17,
	dffe15,
	dffe14,
	pipeline_dffe_16,
	dffe171,
	dffe13,
	pipeline_dffe_15,
	dffe162,
	dffe12,
	pipeline_dffe_14,
	dffe151,
	dffe11,
	pipeline_dffe_13,
	dffe141,
	dffe10,
	pipeline_dffe_12,
	dffe131,
	dffe9,
	pipeline_dffe_11,
	dffe121,
	dffe8,
	pipeline_dffe_10,
	dffe111,
	dffe7,
	pipeline_dffe_9,
	dffe101,
	dffe5,
	dffe6,
	pipeline_dffe_8,
	dffe91,
	pipeline_dffe_7,
	dffe1,
	dffe81,
	dffe2,
	dffe3,
	dffe4,
	pipeline_dffe_6,
	dffe71,
	pipeline_dffe_5,
	dffe61,
	dffe41,
	dffe51,
	pipeline_dffe_4,
	pipeline_dffe_3,
	dffe19,
	dffe21,
	dffe31,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	sin_o_0;
output 	dffe18;
output 	dffe17;
input 	dffe16;
output 	dffe161;
input 	dffe181;
input 	pipeline_dffe_17;
output 	dffe15;
output 	dffe14;
input 	pipeline_dffe_16;
input 	dffe171;
output 	dffe13;
input 	pipeline_dffe_15;
input 	dffe162;
output 	dffe12;
input 	pipeline_dffe_14;
input 	dffe151;
output 	dffe11;
input 	pipeline_dffe_13;
input 	dffe141;
output 	dffe10;
input 	pipeline_dffe_12;
input 	dffe131;
output 	dffe9;
input 	pipeline_dffe_11;
input 	dffe121;
output 	dffe8;
input 	pipeline_dffe_10;
input 	dffe111;
output 	dffe7;
input 	pipeline_dffe_9;
input 	dffe101;
output 	dffe5;
output 	dffe6;
input 	pipeline_dffe_8;
input 	dffe91;
input 	pipeline_dffe_7;
output 	dffe1;
input 	dffe81;
output 	dffe2;
output 	dffe3;
output 	dffe4;
input 	pipeline_dffe_6;
input 	dffe71;
input 	pipeline_dffe_5;
input 	dffe61;
input 	dffe41;
input 	dffe51;
input 	pipeline_dffe_4;
input 	pipeline_dffe_3;
input 	dffe19;
input 	dffe21;
input 	dffe31;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[17]~q ;
wire \xordvalue[14]~q ;
wire \Add0~1_sumout ;
wire \a[16]~q ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \a[15]~q ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \a[14]~q ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \a[13]~q ;
wire \xordvalue[13]~q ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \a[12]~q ;
wire \xordvalue[12]~q ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \a[11]~q ;
wire \xordvalue[11]~q ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \a[10]~q ;
wire \xordvalue[10]~q ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \a[9]~q ;
wire \xordvalue[9]~q ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \a[8]~q ;
wire \xordvalue[8]~q ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \a[7]~q ;
wire \xordvalue[7]~q ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \a[6]~q ;
wire \xordvalue[6]~q ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \a[5]~q ;
wire \xordvalue[5]~q ;
wire \a[4]~q ;
wire \xordvalue[4]~q ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~51 ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~55 ;
wire \a[3]~q ;
wire \xordvalue[3]~q ;
wire \a[0]~q ;
wire \xordvalue[0]~q ;
wire \a[1]~q ;
wire \xordvalue[1]~q ;
wire \a[2]~q ;
wire \xordvalue[2]~q ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~59 ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~63 ;
wire \Add0~65_sumout ;
wire \Add0~66 ;
wire \Add0~67 ;
wire \Add0~69_sumout ;
wire \Add0~70 ;
wire \Add0~71 ;
wire \xordvalue~0_combout ;
wire \xordvalue~1_combout ;
wire \xordvalue~2_combout ;
wire \xordvalue~3_combout ;
wire \xordvalue~4_combout ;
wire \xordvalue~5_combout ;
wire \xordvalue~6_combout ;
wire \xordvalue~7_combout ;
wire \xordvalue~8_combout ;
wire \xordvalue~9_combout ;
wire \xordvalue~10_combout ;
wire \xordvalue~11_combout ;
wire \xordvalue~12_combout ;
wire \xordvalue~13_combout ;
wire \xordvalue~14_combout ;


nco_test_lpm_add_sub_19 u0(
	.a_17(\a[17]~q ),
	.xordvalue_14(\xordvalue[14]~q ),
	.a_16(\a[16]~q ),
	.a_15(\a[15]~q ),
	.a_14(\a[14]~q ),
	.a_13(\a[13]~q ),
	.xordvalue_13(\xordvalue[13]~q ),
	.a_12(\a[12]~q ),
	.xordvalue_12(\xordvalue[12]~q ),
	.a_11(\a[11]~q ),
	.xordvalue_11(\xordvalue[11]~q ),
	.a_10(\a[10]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.a_9(\a[9]~q ),
	.xordvalue_9(\xordvalue[9]~q ),
	.a_8(\a[8]~q ),
	.xordvalue_8(\xordvalue[8]~q ),
	.a_7(\a[7]~q ),
	.xordvalue_7(\xordvalue[7]~q ),
	.a_6(\a[6]~q ),
	.xordvalue_6(\xordvalue[6]~q ),
	.a_5(\a[5]~q ),
	.xordvalue_5(\xordvalue[5]~q ),
	.a_4(\a[4]~q ),
	.xordvalue_4(\xordvalue[4]~q ),
	.a_3(\a[3]~q ),
	.xordvalue_3(\xordvalue[3]~q ),
	.a_0(\a[0]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_1(\a[1]~q ),
	.xordvalue_1(\xordvalue[1]~q ),
	.a_2(\a[2]~q ),
	.xordvalue_2(\xordvalue[2]~q ),
	.dffe18(dffe18),
	.dffe17(dffe17),
	.dffe16(dffe161),
	.dffe15(dffe15),
	.dffe14(dffe14),
	.dffe13(dffe13),
	.dffe12(dffe12),
	.dffe11(dffe11),
	.dffe10(dffe10),
	.dffe9(dffe9),
	.dffe8(dffe8),
	.dffe7(dffe7),
	.dffe5(dffe5),
	.dffe6(dffe6),
	.dffe1(dffe1),
	.dffe2(dffe2),
	.dffe3(dffe3),
	.dffe4(dffe4),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[17] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[17]~q ),
	.prn(vcc));
defparam \a[17] .is_wysiwyg = "true";
defparam \a[17] .power_up = "low";

dffeas \xordvalue[14] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[14]~q ),
	.prn(vcc));
defparam \xordvalue[14] .is_wysiwyg = "true";
defparam \xordvalue[14] .power_up = "low";

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe181),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "on";

dffeas \a[16] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[16]~q ),
	.prn(vcc));
defparam \a[16] .is_wysiwyg = "true";
defparam \a[16] .power_up = "low";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe171),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~5 .shared_arith = "on";

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe162),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~9 .shared_arith = "on";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~13 .shared_arith = "on";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

dffeas \xordvalue[13] (
	.clk(clk),
	.d(\xordvalue~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[13]~q ),
	.prn(vcc));
defparam \xordvalue[13] .is_wysiwyg = "true";
defparam \xordvalue[13] .power_up = "low";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~17 .shared_arith = "on";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

dffeas \xordvalue[12] (
	.clk(clk),
	.d(\xordvalue~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[12]~q ),
	.prn(vcc));
defparam \xordvalue[12] .is_wysiwyg = "true";
defparam \xordvalue[12] .power_up = "low";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "on";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \xordvalue[11] (
	.clk(clk),
	.d(\xordvalue~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[11]~q ),
	.prn(vcc));
defparam \xordvalue[11] .is_wysiwyg = "true";
defparam \xordvalue[11] .power_up = "low";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~25 .shared_arith = "on";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(\xordvalue~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~29 .shared_arith = "on";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \xordvalue[9] (
	.clk(clk),
	.d(\xordvalue~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[9]~q ),
	.prn(vcc));
defparam \xordvalue[9] .is_wysiwyg = "true";
defparam \xordvalue[9] .power_up = "low";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~33 .shared_arith = "on";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \xordvalue[8] (
	.clk(clk),
	.d(\xordvalue~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[8]~q ),
	.prn(vcc));
defparam \xordvalue[8] .is_wysiwyg = "true";
defparam \xordvalue[8] .power_up = "low";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~37 .shared_arith = "on";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \xordvalue[7] (
	.clk(clk),
	.d(\xordvalue~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[7]~q ),
	.prn(vcc));
defparam \xordvalue[7] .is_wysiwyg = "true";
defparam \xordvalue[7] .power_up = "low";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(\Add0~47 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~41 .shared_arith = "on";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \xordvalue[6] (
	.clk(clk),
	.d(\xordvalue~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[6]~q ),
	.prn(vcc));
defparam \xordvalue[6] .is_wysiwyg = "true";
defparam \xordvalue[6] .power_up = "low";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(\Add0~51 ),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout(\Add0~47 ));
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~45 .shared_arith = "on";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \xordvalue[5] (
	.clk(clk),
	.d(\xordvalue~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[5]~q ),
	.prn(vcc));
defparam \xordvalue[5] .is_wysiwyg = "true";
defparam \xordvalue[5] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \xordvalue[4] (
	.clk(clk),
	.d(\xordvalue~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[4]~q ),
	.prn(vcc));
defparam \xordvalue[4] .is_wysiwyg = "true";
defparam \xordvalue[4] .power_up = "low";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(\Add0~55 ),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout(\Add0~51 ));
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~49 .shared_arith = "on";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(\Add0~59 ),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout(\Add0~55 ));
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~53 .shared_arith = "on";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \xordvalue[3] (
	.clk(clk),
	.d(\xordvalue~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[3]~q ),
	.prn(vcc));
defparam \xordvalue[3] .is_wysiwyg = "true";
defparam \xordvalue[3] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \xordvalue[1] (
	.clk(clk),
	.d(\xordvalue~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[1]~q ),
	.prn(vcc));
defparam \xordvalue[1] .is_wysiwyg = "true";
defparam \xordvalue[1] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \xordvalue[2] (
	.clk(clk),
	.d(\xordvalue~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[2]~q ),
	.prn(vcc));
defparam \xordvalue[2] .is_wysiwyg = "true";
defparam \xordvalue[2] .power_up = "low";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~70 ),
	.sharein(\Add0~71 ),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout(\Add0~59 ));
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~57 .shared_arith = "on";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!dffe19),
	.datad(!dffe16),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout(\Add0~63 ));
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add0~61 .shared_arith = "on";

arriav_lcell_comb \Add0~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(\Add0~63 ),
	.combout(),
	.sumout(\Add0~65_sumout ),
	.cout(\Add0~66 ),
	.shareout(\Add0~67 ));
defparam \Add0~65 .extended_lut = "off";
defparam \Add0~65 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~65 .shared_arith = "on";

arriav_lcell_comb \Add0~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~66 ),
	.sharein(\Add0~67 ),
	.combout(),
	.sumout(\Add0~69_sumout ),
	.cout(\Add0~70 ),
	.shareout(\Add0~71 ));
defparam \Add0~69 .extended_lut = "off";
defparam \Add0~69 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~69 .shared_arith = "on";

arriav_lcell_comb \xordvalue~0 (
	.dataa(!pipeline_dffe_17),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

arriav_lcell_comb \xordvalue~1 (
	.dataa(!pipeline_dffe_16),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~1 .extended_lut = "off";
defparam \xordvalue~1 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~1 .shared_arith = "off";

arriav_lcell_comb \xordvalue~2 (
	.dataa(!pipeline_dffe_15),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~2 .extended_lut = "off";
defparam \xordvalue~2 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~2 .shared_arith = "off";

arriav_lcell_comb \xordvalue~3 (
	.dataa(!pipeline_dffe_14),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~3 .extended_lut = "off";
defparam \xordvalue~3 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~3 .shared_arith = "off";

arriav_lcell_comb \xordvalue~4 (
	.dataa(!pipeline_dffe_13),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~4 .extended_lut = "off";
defparam \xordvalue~4 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~4 .shared_arith = "off";

arriav_lcell_comb \xordvalue~5 (
	.dataa(!pipeline_dffe_12),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~5 .extended_lut = "off";
defparam \xordvalue~5 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~5 .shared_arith = "off";

arriav_lcell_comb \xordvalue~6 (
	.dataa(!pipeline_dffe_11),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~6 .extended_lut = "off";
defparam \xordvalue~6 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~6 .shared_arith = "off";

arriav_lcell_comb \xordvalue~7 (
	.dataa(!pipeline_dffe_10),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~7 .extended_lut = "off";
defparam \xordvalue~7 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~7 .shared_arith = "off";

arriav_lcell_comb \xordvalue~8 (
	.dataa(!pipeline_dffe_9),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~8 .extended_lut = "off";
defparam \xordvalue~8 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~8 .shared_arith = "off";

arriav_lcell_comb \xordvalue~9 (
	.dataa(!pipeline_dffe_8),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~9 .extended_lut = "off";
defparam \xordvalue~9 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~9 .shared_arith = "off";

arriav_lcell_comb \xordvalue~10 (
	.dataa(!pipeline_dffe_7),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~10 .extended_lut = "off";
defparam \xordvalue~10 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~10 .shared_arith = "off";

arriav_lcell_comb \xordvalue~11 (
	.dataa(!pipeline_dffe_6),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~11 .extended_lut = "off";
defparam \xordvalue~11 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~11 .shared_arith = "off";

arriav_lcell_comb \xordvalue~12 (
	.dataa(!pipeline_dffe_3),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~12 .extended_lut = "off";
defparam \xordvalue~12 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~12 .shared_arith = "off";

arriav_lcell_comb \xordvalue~13 (
	.dataa(!pipeline_dffe_4),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~13 .extended_lut = "off";
defparam \xordvalue~13 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~13 .shared_arith = "off";

arriav_lcell_comb \xordvalue~14 (
	.dataa(!pipeline_dffe_5),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~14 .extended_lut = "off";
defparam \xordvalue~14 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~14 .shared_arith = "off";

endmodule

module nco_test_lpm_add_sub_19 (
	a_17,
	xordvalue_14,
	a_16,
	a_15,
	a_14,
	a_13,
	xordvalue_13,
	a_12,
	xordvalue_12,
	a_11,
	xordvalue_11,
	a_10,
	xordvalue_10,
	a_9,
	xordvalue_9,
	a_8,
	xordvalue_8,
	a_7,
	xordvalue_7,
	a_6,
	xordvalue_6,
	a_5,
	xordvalue_5,
	a_4,
	xordvalue_4,
	a_3,
	xordvalue_3,
	a_0,
	xordvalue_0,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	dffe18,
	dffe17,
	dffe16,
	dffe15,
	dffe14,
	dffe13,
	dffe12,
	dffe11,
	dffe10,
	dffe9,
	dffe8,
	dffe7,
	dffe5,
	dffe6,
	dffe1,
	dffe2,
	dffe3,
	dffe4,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_14;
input 	a_16;
input 	a_15;
input 	a_14;
input 	a_13;
input 	xordvalue_13;
input 	a_12;
input 	xordvalue_12;
input 	a_11;
input 	xordvalue_11;
input 	a_10;
input 	xordvalue_10;
input 	a_9;
input 	xordvalue_9;
input 	a_8;
input 	xordvalue_8;
input 	a_7;
input 	xordvalue_7;
input 	a_6;
input 	xordvalue_6;
input 	a_5;
input 	xordvalue_5;
input 	a_4;
input 	xordvalue_4;
input 	a_3;
input 	xordvalue_3;
input 	a_0;
input 	xordvalue_0;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
output 	dffe18;
output 	dffe17;
output 	dffe16;
output 	dffe15;
output 	dffe14;
output 	dffe13;
output 	dffe12;
output 	dffe11;
output 	dffe10;
output 	dffe9;
output 	dffe8;
output 	dffe7;
output 	dffe5;
output 	dffe6;
output 	dffe1;
output 	dffe2;
output 	dffe3;
output 	dffe4;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_add_sub_jdg auto_generated(
	.a_17(a_17),
	.xordvalue_14(xordvalue_14),
	.a_16(a_16),
	.a_15(a_15),
	.a_14(a_14),
	.a_13(a_13),
	.xordvalue_13(xordvalue_13),
	.a_12(a_12),
	.xordvalue_12(xordvalue_12),
	.a_11(a_11),
	.xordvalue_11(xordvalue_11),
	.a_10(a_10),
	.xordvalue_10(xordvalue_10),
	.a_9(a_9),
	.xordvalue_9(xordvalue_9),
	.a_8(a_8),
	.xordvalue_8(xordvalue_8),
	.a_7(a_7),
	.xordvalue_7(xordvalue_7),
	.a_6(a_6),
	.xordvalue_6(xordvalue_6),
	.a_5(a_5),
	.xordvalue_5(xordvalue_5),
	.a_4(a_4),
	.xordvalue_4(xordvalue_4),
	.a_3(a_3),
	.xordvalue_3(xordvalue_3),
	.a_0(a_0),
	.xordvalue_0(xordvalue_0),
	.a_1(a_1),
	.xordvalue_1(xordvalue_1),
	.a_2(a_2),
	.xordvalue_2(xordvalue_2),
	.dffe181(dffe18),
	.dffe171(dffe17),
	.dffe161(dffe16),
	.dffe151(dffe15),
	.dffe141(dffe14),
	.dffe131(dffe13),
	.dffe121(dffe12),
	.dffe111(dffe11),
	.dffe101(dffe10),
	.dffe91(dffe9),
	.dffe81(dffe8),
	.dffe71(dffe7),
	.dffe51(dffe5),
	.dffe61(dffe6),
	.dffe19(dffe1),
	.dffe21(dffe2),
	.dffe31(dffe3),
	.dffe41(dffe4),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module nco_test_add_sub_jdg (
	a_17,
	xordvalue_14,
	a_16,
	a_15,
	a_14,
	a_13,
	xordvalue_13,
	a_12,
	xordvalue_12,
	a_11,
	xordvalue_11,
	a_10,
	xordvalue_10,
	a_9,
	xordvalue_9,
	a_8,
	xordvalue_8,
	a_7,
	xordvalue_7,
	a_6,
	xordvalue_6,
	a_5,
	xordvalue_5,
	a_4,
	xordvalue_4,
	a_3,
	xordvalue_3,
	a_0,
	xordvalue_0,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	dffe181,
	dffe171,
	dffe161,
	dffe151,
	dffe141,
	dffe131,
	dffe121,
	dffe111,
	dffe101,
	dffe91,
	dffe81,
	dffe71,
	dffe51,
	dffe61,
	dffe19,
	dffe21,
	dffe31,
	dffe41,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_14;
input 	a_16;
input 	a_15;
input 	a_14;
input 	a_13;
input 	xordvalue_13;
input 	a_12;
input 	xordvalue_12;
input 	a_11;
input 	xordvalue_11;
input 	a_10;
input 	xordvalue_10;
input 	a_9;
input 	xordvalue_9;
input 	a_8;
input 	xordvalue_8;
input 	a_7;
input 	xordvalue_7;
input 	a_6;
input 	xordvalue_6;
input 	a_5;
input 	xordvalue_5;
input 	a_4;
input 	xordvalue_4;
input 	a_3;
input 	xordvalue_3;
input 	a_0;
input 	xordvalue_0;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
output 	dffe181;
output 	dffe171;
output 	dffe161;
output 	dffe151;
output 	dffe141;
output 	dffe131;
output 	dffe121;
output 	dffe111;
output 	dffe101;
output 	dffe91;
output 	dffe81;
output 	dffe71;
output 	dffe51;
output 	dffe61;
output 	dffe19;
output 	dffe21;
output 	dffe31;
output 	dffe41;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~COUT ;
wire \add_sub_cella[12]~COUT ;
wire \add_sub_cella[13]~COUT ;
wire \add_sub_cella[14]~COUT ;
wire \add_sub_cella[15]~COUT ;
wire \add_sub_cella[16]~COUT ;
wire \add_sub_cella[17]~sumout ;
wire \add_sub_cella[16]~sumout ;
wire \add_sub_cella[15]~sumout ;
wire \add_sub_cella[14]~sumout ;
wire \add_sub_cella[13]~sumout ;
wire \add_sub_cella[12]~sumout ;
wire \add_sub_cella[11]~sumout ;
wire \add_sub_cella[10]~sumout ;
wire \add_sub_cella[9]~sumout ;
wire \add_sub_cella[8]~sumout ;
wire \add_sub_cella[7]~sumout ;
wire \add_sub_cella[6]~sumout ;
wire \add_sub_cella[4]~sumout ;
wire \add_sub_cella[5]~sumout ;
wire \add_sub_cella[0]~sumout ;
wire \add_sub_cella[1]~sumout ;
wire \add_sub_cella[2]~sumout ;
wire \add_sub_cella[3]~sumout ;


dffeas dffe18(
	.clk(clock),
	.d(\add_sub_cella[17]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe181),
	.prn(vcc));
defparam dffe18.is_wysiwyg = "true";
defparam dffe18.power_up = "low";

dffeas dffe17(
	.clk(clock),
	.d(\add_sub_cella[16]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe171),
	.prn(vcc));
defparam dffe17.is_wysiwyg = "true";
defparam dffe17.power_up = "low";

dffeas dffe16(
	.clk(clock),
	.d(\add_sub_cella[15]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe161),
	.prn(vcc));
defparam dffe16.is_wysiwyg = "true";
defparam dffe16.power_up = "low";

dffeas dffe15(
	.clk(clock),
	.d(\add_sub_cella[14]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe151),
	.prn(vcc));
defparam dffe15.is_wysiwyg = "true";
defparam dffe15.power_up = "low";

dffeas dffe14(
	.clk(clock),
	.d(\add_sub_cella[13]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe141),
	.prn(vcc));
defparam dffe14.is_wysiwyg = "true";
defparam dffe14.power_up = "low";

dffeas dffe13(
	.clk(clock),
	.d(\add_sub_cella[12]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe131),
	.prn(vcc));
defparam dffe13.is_wysiwyg = "true";
defparam dffe13.power_up = "low";

dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe19),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

arriav_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_1),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_2),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_3),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_4),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_5),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_6),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_7),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_8),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_9),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_11),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(\add_sub_cella[11]~COUT ),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[12] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_12),
	.datag(gnd),
	.cin(\add_sub_cella[11]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[12]~sumout ),
	.cout(\add_sub_cella[12]~COUT ),
	.shareout());
defparam \add_sub_cella[12] .extended_lut = "off";
defparam \add_sub_cella[12] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[12] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[13] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_13),
	.datag(gnd),
	.cin(\add_sub_cella[12]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[13]~sumout ),
	.cout(\add_sub_cella[13]~COUT ),
	.shareout());
defparam \add_sub_cella[13] .extended_lut = "off";
defparam \add_sub_cella[13] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[13] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[14] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_14),
	.datag(gnd),
	.cin(\add_sub_cella[13]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[14]~sumout ),
	.cout(\add_sub_cella[14]~COUT ),
	.shareout());
defparam \add_sub_cella[14] .extended_lut = "off";
defparam \add_sub_cella[14] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[14] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[15] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_14),
	.datag(gnd),
	.cin(\add_sub_cella[14]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[15]~sumout ),
	.cout(\add_sub_cella[15]~COUT ),
	.shareout());
defparam \add_sub_cella[15] .extended_lut = "off";
defparam \add_sub_cella[15] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[15] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[16] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_16),
	.datae(gnd),
	.dataf(!xordvalue_14),
	.datag(gnd),
	.cin(\add_sub_cella[15]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[16]~sumout ),
	.cout(\add_sub_cella[16]~COUT ),
	.shareout());
defparam \add_sub_cella[16] .extended_lut = "off";
defparam \add_sub_cella[16] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[16] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[17] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_17),
	.datae(gnd),
	.dataf(!xordvalue_14),
	.datag(gnd),
	.cin(\add_sub_cella[16]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[17]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[17] .extended_lut = "off";
defparam \add_sub_cella[17] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[17] .shared_arith = "off";

endmodule

module nco_test_cordic_sxor_1p_lpm_1 (
	sin_o_0,
	dffe18,
	dffe17,
	dffe16,
	pipeline_dffe_17,
	dffe161,
	dffe181,
	dffe15,
	dffe171,
	dffe14,
	pipeline_dffe_16,
	dffe162,
	dffe13,
	pipeline_dffe_15,
	dffe151,
	dffe12,
	pipeline_dffe_14,
	dffe141,
	dffe11,
	pipeline_dffe_13,
	dffe131,
	dffe10,
	pipeline_dffe_12,
	dffe121,
	dffe9,
	pipeline_dffe_11,
	dffe111,
	dffe8,
	pipeline_dffe_10,
	dffe6,
	dffe7,
	dffe101,
	pipeline_dffe_9,
	dffe91,
	dffe1,
	pipeline_dffe_8,
	dffe2,
	dffe3,
	dffe4,
	dffe5,
	dffe81,
	pipeline_dffe_7,
	dffe71,
	pipeline_dffe_6,
	dffe51,
	dffe61,
	pipeline_dffe_4,
	pipeline_dffe_5,
	dffe19,
	dffe21,
	dffe31,
	dffe41,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	sin_o_0;
output 	dffe18;
output 	dffe17;
input 	dffe16;
input 	pipeline_dffe_17;
output 	dffe161;
input 	dffe181;
output 	dffe15;
input 	dffe171;
output 	dffe14;
input 	pipeline_dffe_16;
input 	dffe162;
output 	dffe13;
input 	pipeline_dffe_15;
input 	dffe151;
output 	dffe12;
input 	pipeline_dffe_14;
input 	dffe141;
output 	dffe11;
input 	pipeline_dffe_13;
input 	dffe131;
output 	dffe10;
input 	pipeline_dffe_12;
input 	dffe121;
output 	dffe9;
input 	pipeline_dffe_11;
input 	dffe111;
output 	dffe8;
input 	pipeline_dffe_10;
output 	dffe6;
output 	dffe7;
input 	dffe101;
input 	pipeline_dffe_9;
input 	dffe91;
output 	dffe1;
input 	pipeline_dffe_8;
output 	dffe2;
output 	dffe3;
output 	dffe4;
output 	dffe5;
input 	dffe81;
input 	pipeline_dffe_7;
input 	dffe71;
input 	pipeline_dffe_6;
input 	dffe51;
input 	dffe61;
input 	pipeline_dffe_4;
input 	pipeline_dffe_5;
input 	dffe19;
input 	dffe21;
input 	dffe31;
input 	dffe41;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[17]~q ;
wire \xordvalue[13]~q ;
wire \Add0~1_sumout ;
wire \a[16]~q ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \a[15]~q ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \a[14]~q ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \a[13]~q ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \a[12]~q ;
wire \xordvalue[12]~q ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \a[11]~q ;
wire \xordvalue[11]~q ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \a[10]~q ;
wire \xordvalue[10]~q ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \a[9]~q ;
wire \xordvalue[9]~q ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \a[8]~q ;
wire \xordvalue[8]~q ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \a[7]~q ;
wire \xordvalue[7]~q ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \a[6]~q ;
wire \xordvalue[6]~q ;
wire \a[5]~q ;
wire \xordvalue[5]~q ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~51 ;
wire \a[4]~q ;
wire \xordvalue[4]~q ;
wire \a[0]~q ;
wire \xordvalue[0]~q ;
wire \a[1]~q ;
wire \xordvalue[1]~q ;
wire \a[2]~q ;
wire \xordvalue[2]~q ;
wire \a[3]~q ;
wire \xordvalue[3]~q ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~55 ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~59 ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~63 ;
wire \Add0~65_sumout ;
wire \Add0~66 ;
wire \Add0~67 ;
wire \Add0~69_sumout ;
wire \Add0~70 ;
wire \Add0~71 ;
wire \xordvalue~0_combout ;
wire \xordvalue~1_combout ;
wire \xordvalue~2_combout ;
wire \xordvalue~3_combout ;
wire \xordvalue~4_combout ;
wire \xordvalue~5_combout ;
wire \xordvalue~6_combout ;
wire \xordvalue~7_combout ;
wire \xordvalue~8_combout ;
wire \xordvalue~9_combout ;
wire \xordvalue~10_combout ;
wire \xordvalue~11_combout ;
wire \xordvalue~12_combout ;
wire \xordvalue~13_combout ;


nco_test_lpm_add_sub_20 u0(
	.a_17(\a[17]~q ),
	.xordvalue_13(\xordvalue[13]~q ),
	.a_16(\a[16]~q ),
	.a_15(\a[15]~q ),
	.a_14(\a[14]~q ),
	.a_13(\a[13]~q ),
	.a_12(\a[12]~q ),
	.xordvalue_12(\xordvalue[12]~q ),
	.a_11(\a[11]~q ),
	.xordvalue_11(\xordvalue[11]~q ),
	.a_10(\a[10]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.a_9(\a[9]~q ),
	.xordvalue_9(\xordvalue[9]~q ),
	.a_8(\a[8]~q ),
	.xordvalue_8(\xordvalue[8]~q ),
	.a_7(\a[7]~q ),
	.xordvalue_7(\xordvalue[7]~q ),
	.a_6(\a[6]~q ),
	.xordvalue_6(\xordvalue[6]~q ),
	.a_5(\a[5]~q ),
	.xordvalue_5(\xordvalue[5]~q ),
	.a_4(\a[4]~q ),
	.xordvalue_4(\xordvalue[4]~q ),
	.a_0(\a[0]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_1(\a[1]~q ),
	.xordvalue_1(\xordvalue[1]~q ),
	.a_2(\a[2]~q ),
	.xordvalue_2(\xordvalue[2]~q ),
	.a_3(\a[3]~q ),
	.xordvalue_3(\xordvalue[3]~q ),
	.dffe18(dffe18),
	.dffe17(dffe17),
	.dffe16(dffe161),
	.dffe15(dffe15),
	.dffe14(dffe14),
	.dffe13(dffe13),
	.dffe12(dffe12),
	.dffe11(dffe11),
	.dffe10(dffe10),
	.dffe9(dffe9),
	.dffe8(dffe8),
	.dffe6(dffe6),
	.dffe7(dffe7),
	.dffe1(dffe1),
	.dffe2(dffe2),
	.dffe3(dffe3),
	.dffe4(dffe4),
	.dffe5(dffe5),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[17] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[17]~q ),
	.prn(vcc));
defparam \a[17] .is_wysiwyg = "true";
defparam \a[17] .power_up = "low";

dffeas \xordvalue[13] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[13]~q ),
	.prn(vcc));
defparam \xordvalue[13] .is_wysiwyg = "true";
defparam \xordvalue[13] .power_up = "low";

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe181),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "on";

dffeas \a[16] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[16]~q ),
	.prn(vcc));
defparam \a[16] .is_wysiwyg = "true";
defparam \a[16] .power_up = "low";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe171),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~5 .shared_arith = "on";

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe162),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~9 .shared_arith = "on";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~13 .shared_arith = "on";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~17 .shared_arith = "on";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

dffeas \xordvalue[12] (
	.clk(clk),
	.d(\xordvalue~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[12]~q ),
	.prn(vcc));
defparam \xordvalue[12] .is_wysiwyg = "true";
defparam \xordvalue[12] .power_up = "low";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "on";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \xordvalue[11] (
	.clk(clk),
	.d(\xordvalue~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[11]~q ),
	.prn(vcc));
defparam \xordvalue[11] .is_wysiwyg = "true";
defparam \xordvalue[11] .power_up = "low";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~25 .shared_arith = "on";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(\xordvalue~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~29 .shared_arith = "on";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \xordvalue[9] (
	.clk(clk),
	.d(\xordvalue~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[9]~q ),
	.prn(vcc));
defparam \xordvalue[9] .is_wysiwyg = "true";
defparam \xordvalue[9] .power_up = "low";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~33 .shared_arith = "on";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \xordvalue[8] (
	.clk(clk),
	.d(\xordvalue~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[8]~q ),
	.prn(vcc));
defparam \xordvalue[8] .is_wysiwyg = "true";
defparam \xordvalue[8] .power_up = "low";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~37 .shared_arith = "on";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \xordvalue[7] (
	.clk(clk),
	.d(\xordvalue~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[7]~q ),
	.prn(vcc));
defparam \xordvalue[7] .is_wysiwyg = "true";
defparam \xordvalue[7] .power_up = "low";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(\Add0~47 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~41 .shared_arith = "on";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \xordvalue[6] (
	.clk(clk),
	.d(\xordvalue~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[6]~q ),
	.prn(vcc));
defparam \xordvalue[6] .is_wysiwyg = "true";
defparam \xordvalue[6] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \xordvalue[5] (
	.clk(clk),
	.d(\xordvalue~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[5]~q ),
	.prn(vcc));
defparam \xordvalue[5] .is_wysiwyg = "true";
defparam \xordvalue[5] .power_up = "low";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(\Add0~51 ),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout(\Add0~47 ));
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~45 .shared_arith = "on";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(\Add0~55 ),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout(\Add0~51 ));
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~49 .shared_arith = "on";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \xordvalue[4] (
	.clk(clk),
	.d(\xordvalue~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[4]~q ),
	.prn(vcc));
defparam \xordvalue[4] .is_wysiwyg = "true";
defparam \xordvalue[4] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \xordvalue[1] (
	.clk(clk),
	.d(\xordvalue~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[1]~q ),
	.prn(vcc));
defparam \xordvalue[1] .is_wysiwyg = "true";
defparam \xordvalue[1] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \xordvalue[2] (
	.clk(clk),
	.d(\xordvalue~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[2]~q ),
	.prn(vcc));
defparam \xordvalue[2] .is_wysiwyg = "true";
defparam \xordvalue[2] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \xordvalue[3] (
	.clk(clk),
	.d(\xordvalue~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[3]~q ),
	.prn(vcc));
defparam \xordvalue[3] .is_wysiwyg = "true";
defparam \xordvalue[3] .power_up = "low";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~70 ),
	.sharein(\Add0~71 ),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout(\Add0~55 ));
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~53 .shared_arith = "on";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!dffe19),
	.datad(!dffe16),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout(\Add0~59 ));
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add0~57 .shared_arith = "on";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(\Add0~59 ),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout(\Add0~63 ));
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~61 .shared_arith = "on";

arriav_lcell_comb \Add0~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(\Add0~63 ),
	.combout(),
	.sumout(\Add0~65_sumout ),
	.cout(\Add0~66 ),
	.shareout(\Add0~67 ));
defparam \Add0~65 .extended_lut = "off";
defparam \Add0~65 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~65 .shared_arith = "on";

arriav_lcell_comb \Add0~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~66 ),
	.sharein(\Add0~67 ),
	.combout(),
	.sumout(\Add0~69_sumout ),
	.cout(\Add0~70 ),
	.shareout(\Add0~71 ));
defparam \Add0~69 .extended_lut = "off";
defparam \Add0~69 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~69 .shared_arith = "on";

arriav_lcell_comb \xordvalue~0 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_17),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

arriav_lcell_comb \xordvalue~1 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~1 .extended_lut = "off";
defparam \xordvalue~1 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~1 .shared_arith = "off";

arriav_lcell_comb \xordvalue~2 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_15),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~2 .extended_lut = "off";
defparam \xordvalue~2 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~2 .shared_arith = "off";

arriav_lcell_comb \xordvalue~3 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_14),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~3 .extended_lut = "off";
defparam \xordvalue~3 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~3 .shared_arith = "off";

arriav_lcell_comb \xordvalue~4 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_13),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~4 .extended_lut = "off";
defparam \xordvalue~4 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~4 .shared_arith = "off";

arriav_lcell_comb \xordvalue~5 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_12),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~5 .extended_lut = "off";
defparam \xordvalue~5 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~5 .shared_arith = "off";

arriav_lcell_comb \xordvalue~6 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_11),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~6 .extended_lut = "off";
defparam \xordvalue~6 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~6 .shared_arith = "off";

arriav_lcell_comb \xordvalue~7 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_10),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~7 .extended_lut = "off";
defparam \xordvalue~7 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~7 .shared_arith = "off";

arriav_lcell_comb \xordvalue~8 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_9),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~8 .extended_lut = "off";
defparam \xordvalue~8 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~8 .shared_arith = "off";

arriav_lcell_comb \xordvalue~9 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_8),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~9 .extended_lut = "off";
defparam \xordvalue~9 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~9 .shared_arith = "off";

arriav_lcell_comb \xordvalue~10 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_4),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~10 .extended_lut = "off";
defparam \xordvalue~10 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~10 .shared_arith = "off";

arriav_lcell_comb \xordvalue~11 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_5),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~11 .extended_lut = "off";
defparam \xordvalue~11 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~11 .shared_arith = "off";

arriav_lcell_comb \xordvalue~12 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_6),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~12 .extended_lut = "off";
defparam \xordvalue~12 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~12 .shared_arith = "off";

arriav_lcell_comb \xordvalue~13 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_7),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~13 .extended_lut = "off";
defparam \xordvalue~13 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~13 .shared_arith = "off";

endmodule

module nco_test_lpm_add_sub_20 (
	a_17,
	xordvalue_13,
	a_16,
	a_15,
	a_14,
	a_13,
	a_12,
	xordvalue_12,
	a_11,
	xordvalue_11,
	a_10,
	xordvalue_10,
	a_9,
	xordvalue_9,
	a_8,
	xordvalue_8,
	a_7,
	xordvalue_7,
	a_6,
	xordvalue_6,
	a_5,
	xordvalue_5,
	a_4,
	xordvalue_4,
	a_0,
	xordvalue_0,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	dffe18,
	dffe17,
	dffe16,
	dffe15,
	dffe14,
	dffe13,
	dffe12,
	dffe11,
	dffe10,
	dffe9,
	dffe8,
	dffe6,
	dffe7,
	dffe1,
	dffe2,
	dffe3,
	dffe4,
	dffe5,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_13;
input 	a_16;
input 	a_15;
input 	a_14;
input 	a_13;
input 	a_12;
input 	xordvalue_12;
input 	a_11;
input 	xordvalue_11;
input 	a_10;
input 	xordvalue_10;
input 	a_9;
input 	xordvalue_9;
input 	a_8;
input 	xordvalue_8;
input 	a_7;
input 	xordvalue_7;
input 	a_6;
input 	xordvalue_6;
input 	a_5;
input 	xordvalue_5;
input 	a_4;
input 	xordvalue_4;
input 	a_0;
input 	xordvalue_0;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
output 	dffe18;
output 	dffe17;
output 	dffe16;
output 	dffe15;
output 	dffe14;
output 	dffe13;
output 	dffe12;
output 	dffe11;
output 	dffe10;
output 	dffe9;
output 	dffe8;
output 	dffe6;
output 	dffe7;
output 	dffe1;
output 	dffe2;
output 	dffe3;
output 	dffe4;
output 	dffe5;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_add_sub_jdg_1 auto_generated(
	.a_17(a_17),
	.xordvalue_13(xordvalue_13),
	.a_16(a_16),
	.a_15(a_15),
	.a_14(a_14),
	.a_13(a_13),
	.a_12(a_12),
	.xordvalue_12(xordvalue_12),
	.a_11(a_11),
	.xordvalue_11(xordvalue_11),
	.a_10(a_10),
	.xordvalue_10(xordvalue_10),
	.a_9(a_9),
	.xordvalue_9(xordvalue_9),
	.a_8(a_8),
	.xordvalue_8(xordvalue_8),
	.a_7(a_7),
	.xordvalue_7(xordvalue_7),
	.a_6(a_6),
	.xordvalue_6(xordvalue_6),
	.a_5(a_5),
	.xordvalue_5(xordvalue_5),
	.a_4(a_4),
	.xordvalue_4(xordvalue_4),
	.a_0(a_0),
	.xordvalue_0(xordvalue_0),
	.a_1(a_1),
	.xordvalue_1(xordvalue_1),
	.a_2(a_2),
	.xordvalue_2(xordvalue_2),
	.a_3(a_3),
	.xordvalue_3(xordvalue_3),
	.dffe181(dffe18),
	.dffe171(dffe17),
	.dffe161(dffe16),
	.dffe151(dffe15),
	.dffe141(dffe14),
	.dffe131(dffe13),
	.dffe121(dffe12),
	.dffe111(dffe11),
	.dffe101(dffe10),
	.dffe91(dffe9),
	.dffe81(dffe8),
	.dffe61(dffe6),
	.dffe71(dffe7),
	.dffe19(dffe1),
	.dffe21(dffe2),
	.dffe31(dffe3),
	.dffe41(dffe4),
	.dffe51(dffe5),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module nco_test_add_sub_jdg_1 (
	a_17,
	xordvalue_13,
	a_16,
	a_15,
	a_14,
	a_13,
	a_12,
	xordvalue_12,
	a_11,
	xordvalue_11,
	a_10,
	xordvalue_10,
	a_9,
	xordvalue_9,
	a_8,
	xordvalue_8,
	a_7,
	xordvalue_7,
	a_6,
	xordvalue_6,
	a_5,
	xordvalue_5,
	a_4,
	xordvalue_4,
	a_0,
	xordvalue_0,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	dffe181,
	dffe171,
	dffe161,
	dffe151,
	dffe141,
	dffe131,
	dffe121,
	dffe111,
	dffe101,
	dffe91,
	dffe81,
	dffe61,
	dffe71,
	dffe19,
	dffe21,
	dffe31,
	dffe41,
	dffe51,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_13;
input 	a_16;
input 	a_15;
input 	a_14;
input 	a_13;
input 	a_12;
input 	xordvalue_12;
input 	a_11;
input 	xordvalue_11;
input 	a_10;
input 	xordvalue_10;
input 	a_9;
input 	xordvalue_9;
input 	a_8;
input 	xordvalue_8;
input 	a_7;
input 	xordvalue_7;
input 	a_6;
input 	xordvalue_6;
input 	a_5;
input 	xordvalue_5;
input 	a_4;
input 	xordvalue_4;
input 	a_0;
input 	xordvalue_0;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
output 	dffe181;
output 	dffe171;
output 	dffe161;
output 	dffe151;
output 	dffe141;
output 	dffe131;
output 	dffe121;
output 	dffe111;
output 	dffe101;
output 	dffe91;
output 	dffe81;
output 	dffe61;
output 	dffe71;
output 	dffe19;
output 	dffe21;
output 	dffe31;
output 	dffe41;
output 	dffe51;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~COUT ;
wire \add_sub_cella[12]~COUT ;
wire \add_sub_cella[13]~COUT ;
wire \add_sub_cella[14]~COUT ;
wire \add_sub_cella[15]~COUT ;
wire \add_sub_cella[16]~COUT ;
wire \add_sub_cella[17]~sumout ;
wire \add_sub_cella[16]~sumout ;
wire \add_sub_cella[15]~sumout ;
wire \add_sub_cella[14]~sumout ;
wire \add_sub_cella[13]~sumout ;
wire \add_sub_cella[12]~sumout ;
wire \add_sub_cella[11]~sumout ;
wire \add_sub_cella[10]~sumout ;
wire \add_sub_cella[9]~sumout ;
wire \add_sub_cella[8]~sumout ;
wire \add_sub_cella[7]~sumout ;
wire \add_sub_cella[5]~sumout ;
wire \add_sub_cella[6]~sumout ;
wire \add_sub_cella[0]~sumout ;
wire \add_sub_cella[1]~sumout ;
wire \add_sub_cella[2]~sumout ;
wire \add_sub_cella[3]~sumout ;
wire \add_sub_cella[4]~sumout ;


dffeas dffe18(
	.clk(clock),
	.d(\add_sub_cella[17]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe181),
	.prn(vcc));
defparam dffe18.is_wysiwyg = "true";
defparam dffe18.power_up = "low";

dffeas dffe17(
	.clk(clock),
	.d(\add_sub_cella[16]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe171),
	.prn(vcc));
defparam dffe17.is_wysiwyg = "true";
defparam dffe17.power_up = "low";

dffeas dffe16(
	.clk(clock),
	.d(\add_sub_cella[15]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe161),
	.prn(vcc));
defparam dffe16.is_wysiwyg = "true";
defparam dffe16.power_up = "low";

dffeas dffe15(
	.clk(clock),
	.d(\add_sub_cella[14]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe151),
	.prn(vcc));
defparam dffe15.is_wysiwyg = "true";
defparam dffe15.power_up = "low";

dffeas dffe14(
	.clk(clock),
	.d(\add_sub_cella[13]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe141),
	.prn(vcc));
defparam dffe14.is_wysiwyg = "true";
defparam dffe14.power_up = "low";

dffeas dffe13(
	.clk(clock),
	.d(\add_sub_cella[12]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe131),
	.prn(vcc));
defparam dffe13.is_wysiwyg = "true";
defparam dffe13.power_up = "low";

dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe19),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

arriav_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_1),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_2),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_3),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_4),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_5),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_6),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_7),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_8),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_9),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_11),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(\add_sub_cella[11]~COUT ),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[12] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_12),
	.datag(gnd),
	.cin(\add_sub_cella[11]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[12]~sumout ),
	.cout(\add_sub_cella[12]~COUT ),
	.shareout());
defparam \add_sub_cella[12] .extended_lut = "off";
defparam \add_sub_cella[12] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[12] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[13] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_13),
	.datag(gnd),
	.cin(\add_sub_cella[12]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[13]~sumout ),
	.cout(\add_sub_cella[13]~COUT ),
	.shareout());
defparam \add_sub_cella[13] .extended_lut = "off";
defparam \add_sub_cella[13] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[13] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[14] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_13),
	.datag(gnd),
	.cin(\add_sub_cella[13]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[14]~sumout ),
	.cout(\add_sub_cella[14]~COUT ),
	.shareout());
defparam \add_sub_cella[14] .extended_lut = "off";
defparam \add_sub_cella[14] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[14] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[15] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_13),
	.datag(gnd),
	.cin(\add_sub_cella[14]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[15]~sumout ),
	.cout(\add_sub_cella[15]~COUT ),
	.shareout());
defparam \add_sub_cella[15] .extended_lut = "off";
defparam \add_sub_cella[15] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[15] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[16] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_16),
	.datae(gnd),
	.dataf(!xordvalue_13),
	.datag(gnd),
	.cin(\add_sub_cella[15]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[16]~sumout ),
	.cout(\add_sub_cella[16]~COUT ),
	.shareout());
defparam \add_sub_cella[16] .extended_lut = "off";
defparam \add_sub_cella[16] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[16] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[17] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_17),
	.datae(gnd),
	.dataf(!xordvalue_13),
	.datag(gnd),
	.cin(\add_sub_cella[16]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[17]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[17] .extended_lut = "off";
defparam \add_sub_cella[17] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[17] .shared_arith = "off";

endmodule

module nco_test_cordic_sxor_1p_lpm_2 (
	sin_o_0,
	dffe18,
	dffe17,
	dffe16,
	dffe161,
	dffe181,
	pipeline_dffe_17,
	dffe15,
	dffe14,
	pipeline_dffe_16,
	dffe171,
	dffe13,
	pipeline_dffe_15,
	dffe162,
	dffe12,
	pipeline_dffe_14,
	dffe151,
	dffe11,
	pipeline_dffe_13,
	dffe141,
	dffe10,
	pipeline_dffe_12,
	dffe131,
	dffe9,
	pipeline_dffe_11,
	dffe121,
	dffe7,
	dffe8,
	pipeline_dffe_10,
	dffe111,
	pipeline_dffe_9,
	dffe1,
	dffe101,
	dffe2,
	dffe3,
	dffe4,
	dffe5,
	dffe6,
	pipeline_dffe_8,
	dffe91,
	pipeline_dffe_7,
	dffe81,
	dffe61,
	dffe71,
	pipeline_dffe_6,
	pipeline_dffe_5,
	dffe19,
	dffe21,
	dffe31,
	dffe41,
	dffe51,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	sin_o_0;
output 	dffe18;
output 	dffe17;
input 	dffe16;
output 	dffe161;
input 	dffe181;
input 	pipeline_dffe_17;
output 	dffe15;
output 	dffe14;
input 	pipeline_dffe_16;
input 	dffe171;
output 	dffe13;
input 	pipeline_dffe_15;
input 	dffe162;
output 	dffe12;
input 	pipeline_dffe_14;
input 	dffe151;
output 	dffe11;
input 	pipeline_dffe_13;
input 	dffe141;
output 	dffe10;
input 	pipeline_dffe_12;
input 	dffe131;
output 	dffe9;
input 	pipeline_dffe_11;
input 	dffe121;
output 	dffe7;
output 	dffe8;
input 	pipeline_dffe_10;
input 	dffe111;
input 	pipeline_dffe_9;
output 	dffe1;
input 	dffe101;
output 	dffe2;
output 	dffe3;
output 	dffe4;
output 	dffe5;
output 	dffe6;
input 	pipeline_dffe_8;
input 	dffe91;
input 	pipeline_dffe_7;
input 	dffe81;
input 	dffe61;
input 	dffe71;
input 	pipeline_dffe_6;
input 	pipeline_dffe_5;
input 	dffe19;
input 	dffe21;
input 	dffe31;
input 	dffe41;
input 	dffe51;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[17]~q ;
wire \xordvalue[12]~q ;
wire \Add0~1_sumout ;
wire \a[16]~q ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \a[15]~q ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \a[14]~q ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \a[13]~q ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \a[12]~q ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \a[11]~q ;
wire \xordvalue[11]~q ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \a[10]~q ;
wire \xordvalue[10]~q ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \a[9]~q ;
wire \xordvalue[9]~q ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \a[8]~q ;
wire \xordvalue[8]~q ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \a[7]~q ;
wire \xordvalue[7]~q ;
wire \a[6]~q ;
wire \xordvalue[6]~q ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \a[5]~q ;
wire \xordvalue[5]~q ;
wire \a[0]~q ;
wire \xordvalue[0]~q ;
wire \a[1]~q ;
wire \xordvalue[1]~q ;
wire \a[2]~q ;
wire \xordvalue[2]~q ;
wire \a[3]~q ;
wire \xordvalue[3]~q ;
wire \a[4]~q ;
wire \xordvalue[4]~q ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~51 ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~55 ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~59 ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~63 ;
wire \Add0~65_sumout ;
wire \Add0~66 ;
wire \Add0~67 ;
wire \Add0~69_sumout ;
wire \Add0~70 ;
wire \Add0~71 ;
wire \xordvalue~0_combout ;
wire \xordvalue~1_combout ;
wire \xordvalue~2_combout ;
wire \xordvalue~3_combout ;
wire \xordvalue~4_combout ;
wire \xordvalue~5_combout ;
wire \xordvalue~6_combout ;
wire \xordvalue~7_combout ;
wire \xordvalue~8_combout ;
wire \xordvalue~9_combout ;
wire \xordvalue~10_combout ;
wire \xordvalue~11_combout ;
wire \xordvalue~12_combout ;


nco_test_lpm_add_sub_21 u0(
	.a_17(\a[17]~q ),
	.xordvalue_12(\xordvalue[12]~q ),
	.a_16(\a[16]~q ),
	.a_15(\a[15]~q ),
	.a_14(\a[14]~q ),
	.a_13(\a[13]~q ),
	.a_12(\a[12]~q ),
	.a_11(\a[11]~q ),
	.xordvalue_11(\xordvalue[11]~q ),
	.a_10(\a[10]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.a_9(\a[9]~q ),
	.xordvalue_9(\xordvalue[9]~q ),
	.a_8(\a[8]~q ),
	.xordvalue_8(\xordvalue[8]~q ),
	.a_7(\a[7]~q ),
	.xordvalue_7(\xordvalue[7]~q ),
	.a_6(\a[6]~q ),
	.xordvalue_6(\xordvalue[6]~q ),
	.a_5(\a[5]~q ),
	.xordvalue_5(\xordvalue[5]~q ),
	.a_0(\a[0]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_1(\a[1]~q ),
	.xordvalue_1(\xordvalue[1]~q ),
	.a_2(\a[2]~q ),
	.xordvalue_2(\xordvalue[2]~q ),
	.a_3(\a[3]~q ),
	.xordvalue_3(\xordvalue[3]~q ),
	.a_4(\a[4]~q ),
	.xordvalue_4(\xordvalue[4]~q ),
	.dffe18(dffe18),
	.dffe17(dffe17),
	.dffe16(dffe161),
	.dffe15(dffe15),
	.dffe14(dffe14),
	.dffe13(dffe13),
	.dffe12(dffe12),
	.dffe11(dffe11),
	.dffe10(dffe10),
	.dffe9(dffe9),
	.dffe7(dffe7),
	.dffe8(dffe8),
	.dffe1(dffe1),
	.dffe2(dffe2),
	.dffe3(dffe3),
	.dffe4(dffe4),
	.dffe5(dffe5),
	.dffe6(dffe6),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[17] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[17]~q ),
	.prn(vcc));
defparam \a[17] .is_wysiwyg = "true";
defparam \a[17] .power_up = "low";

dffeas \xordvalue[12] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[12]~q ),
	.prn(vcc));
defparam \xordvalue[12] .is_wysiwyg = "true";
defparam \xordvalue[12] .power_up = "low";

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe181),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "on";

dffeas \a[16] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[16]~q ),
	.prn(vcc));
defparam \a[16] .is_wysiwyg = "true";
defparam \a[16] .power_up = "low";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe171),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~5 .shared_arith = "on";

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe162),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~9 .shared_arith = "on";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~13 .shared_arith = "on";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~17 .shared_arith = "on";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "on";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \xordvalue[11] (
	.clk(clk),
	.d(\xordvalue~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[11]~q ),
	.prn(vcc));
defparam \xordvalue[11] .is_wysiwyg = "true";
defparam \xordvalue[11] .power_up = "low";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~25 .shared_arith = "on";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(\xordvalue~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~29 .shared_arith = "on";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \xordvalue[9] (
	.clk(clk),
	.d(\xordvalue~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[9]~q ),
	.prn(vcc));
defparam \xordvalue[9] .is_wysiwyg = "true";
defparam \xordvalue[9] .power_up = "low";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~33 .shared_arith = "on";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \xordvalue[8] (
	.clk(clk),
	.d(\xordvalue~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[8]~q ),
	.prn(vcc));
defparam \xordvalue[8] .is_wysiwyg = "true";
defparam \xordvalue[8] .power_up = "low";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~37 .shared_arith = "on";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \xordvalue[7] (
	.clk(clk),
	.d(\xordvalue~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[7]~q ),
	.prn(vcc));
defparam \xordvalue[7] .is_wysiwyg = "true";
defparam \xordvalue[7] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \xordvalue[6] (
	.clk(clk),
	.d(\xordvalue~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[6]~q ),
	.prn(vcc));
defparam \xordvalue[6] .is_wysiwyg = "true";
defparam \xordvalue[6] .power_up = "low";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(\Add0~47 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~41 .shared_arith = "on";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(\Add0~51 ),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout(\Add0~47 ));
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~45 .shared_arith = "on";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \xordvalue[5] (
	.clk(clk),
	.d(\xordvalue~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[5]~q ),
	.prn(vcc));
defparam \xordvalue[5] .is_wysiwyg = "true";
defparam \xordvalue[5] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \xordvalue[1] (
	.clk(clk),
	.d(\xordvalue~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[1]~q ),
	.prn(vcc));
defparam \xordvalue[1] .is_wysiwyg = "true";
defparam \xordvalue[1] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \xordvalue[2] (
	.clk(clk),
	.d(\xordvalue~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[2]~q ),
	.prn(vcc));
defparam \xordvalue[2] .is_wysiwyg = "true";
defparam \xordvalue[2] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \xordvalue[3] (
	.clk(clk),
	.d(\xordvalue~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[3]~q ),
	.prn(vcc));
defparam \xordvalue[3] .is_wysiwyg = "true";
defparam \xordvalue[3] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \xordvalue[4] (
	.clk(clk),
	.d(\xordvalue~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[4]~q ),
	.prn(vcc));
defparam \xordvalue[4] .is_wysiwyg = "true";
defparam \xordvalue[4] .power_up = "low";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~70 ),
	.sharein(\Add0~71 ),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout(\Add0~51 ));
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~49 .shared_arith = "on";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!dffe19),
	.datad(!dffe16),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout(\Add0~55 ));
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add0~53 .shared_arith = "on";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(\Add0~55 ),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout(\Add0~59 ));
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~57 .shared_arith = "on";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(\Add0~59 ),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout(\Add0~63 ));
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~61 .shared_arith = "on";

arriav_lcell_comb \Add0~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(\Add0~63 ),
	.combout(),
	.sumout(\Add0~65_sumout ),
	.cout(\Add0~66 ),
	.shareout(\Add0~67 ));
defparam \Add0~65 .extended_lut = "off";
defparam \Add0~65 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~65 .shared_arith = "on";

arriav_lcell_comb \Add0~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~66 ),
	.sharein(\Add0~67 ),
	.combout(),
	.sumout(\Add0~69_sumout ),
	.cout(\Add0~70 ),
	.shareout(\Add0~71 ));
defparam \Add0~69 .extended_lut = "off";
defparam \Add0~69 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~69 .shared_arith = "on";

arriav_lcell_comb \xordvalue~0 (
	.dataa(!pipeline_dffe_17),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

arriav_lcell_comb \xordvalue~1 (
	.dataa(!pipeline_dffe_16),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~1 .extended_lut = "off";
defparam \xordvalue~1 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~1 .shared_arith = "off";

arriav_lcell_comb \xordvalue~2 (
	.dataa(!pipeline_dffe_15),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~2 .extended_lut = "off";
defparam \xordvalue~2 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~2 .shared_arith = "off";

arriav_lcell_comb \xordvalue~3 (
	.dataa(!pipeline_dffe_14),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~3 .extended_lut = "off";
defparam \xordvalue~3 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~3 .shared_arith = "off";

arriav_lcell_comb \xordvalue~4 (
	.dataa(!pipeline_dffe_13),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~4 .extended_lut = "off";
defparam \xordvalue~4 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~4 .shared_arith = "off";

arriav_lcell_comb \xordvalue~5 (
	.dataa(!pipeline_dffe_12),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~5 .extended_lut = "off";
defparam \xordvalue~5 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~5 .shared_arith = "off";

arriav_lcell_comb \xordvalue~6 (
	.dataa(!pipeline_dffe_11),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~6 .extended_lut = "off";
defparam \xordvalue~6 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~6 .shared_arith = "off";

arriav_lcell_comb \xordvalue~7 (
	.dataa(!pipeline_dffe_10),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~7 .extended_lut = "off";
defparam \xordvalue~7 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~7 .shared_arith = "off";

arriav_lcell_comb \xordvalue~8 (
	.dataa(!pipeline_dffe_5),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~8 .extended_lut = "off";
defparam \xordvalue~8 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~8 .shared_arith = "off";

arriav_lcell_comb \xordvalue~9 (
	.dataa(!pipeline_dffe_6),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~9 .extended_lut = "off";
defparam \xordvalue~9 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~9 .shared_arith = "off";

arriav_lcell_comb \xordvalue~10 (
	.dataa(!pipeline_dffe_7),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~10 .extended_lut = "off";
defparam \xordvalue~10 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~10 .shared_arith = "off";

arriav_lcell_comb \xordvalue~11 (
	.dataa(!pipeline_dffe_8),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~11 .extended_lut = "off";
defparam \xordvalue~11 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~11 .shared_arith = "off";

arriav_lcell_comb \xordvalue~12 (
	.dataa(!pipeline_dffe_9),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~12 .extended_lut = "off";
defparam \xordvalue~12 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~12 .shared_arith = "off";

endmodule

module nco_test_lpm_add_sub_21 (
	a_17,
	xordvalue_12,
	a_16,
	a_15,
	a_14,
	a_13,
	a_12,
	a_11,
	xordvalue_11,
	a_10,
	xordvalue_10,
	a_9,
	xordvalue_9,
	a_8,
	xordvalue_8,
	a_7,
	xordvalue_7,
	a_6,
	xordvalue_6,
	a_5,
	xordvalue_5,
	a_0,
	xordvalue_0,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	a_4,
	xordvalue_4,
	dffe18,
	dffe17,
	dffe16,
	dffe15,
	dffe14,
	dffe13,
	dffe12,
	dffe11,
	dffe10,
	dffe9,
	dffe7,
	dffe8,
	dffe1,
	dffe2,
	dffe3,
	dffe4,
	dffe5,
	dffe6,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_12;
input 	a_16;
input 	a_15;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	xordvalue_11;
input 	a_10;
input 	xordvalue_10;
input 	a_9;
input 	xordvalue_9;
input 	a_8;
input 	xordvalue_8;
input 	a_7;
input 	xordvalue_7;
input 	a_6;
input 	xordvalue_6;
input 	a_5;
input 	xordvalue_5;
input 	a_0;
input 	xordvalue_0;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
input 	a_4;
input 	xordvalue_4;
output 	dffe18;
output 	dffe17;
output 	dffe16;
output 	dffe15;
output 	dffe14;
output 	dffe13;
output 	dffe12;
output 	dffe11;
output 	dffe10;
output 	dffe9;
output 	dffe7;
output 	dffe8;
output 	dffe1;
output 	dffe2;
output 	dffe3;
output 	dffe4;
output 	dffe5;
output 	dffe6;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_add_sub_jdg_2 auto_generated(
	.a_17(a_17),
	.xordvalue_12(xordvalue_12),
	.a_16(a_16),
	.a_15(a_15),
	.a_14(a_14),
	.a_13(a_13),
	.a_12(a_12),
	.a_11(a_11),
	.xordvalue_11(xordvalue_11),
	.a_10(a_10),
	.xordvalue_10(xordvalue_10),
	.a_9(a_9),
	.xordvalue_9(xordvalue_9),
	.a_8(a_8),
	.xordvalue_8(xordvalue_8),
	.a_7(a_7),
	.xordvalue_7(xordvalue_7),
	.a_6(a_6),
	.xordvalue_6(xordvalue_6),
	.a_5(a_5),
	.xordvalue_5(xordvalue_5),
	.a_0(a_0),
	.xordvalue_0(xordvalue_0),
	.a_1(a_1),
	.xordvalue_1(xordvalue_1),
	.a_2(a_2),
	.xordvalue_2(xordvalue_2),
	.a_3(a_3),
	.xordvalue_3(xordvalue_3),
	.a_4(a_4),
	.xordvalue_4(xordvalue_4),
	.dffe181(dffe18),
	.dffe171(dffe17),
	.dffe161(dffe16),
	.dffe151(dffe15),
	.dffe141(dffe14),
	.dffe131(dffe13),
	.dffe121(dffe12),
	.dffe111(dffe11),
	.dffe101(dffe10),
	.dffe91(dffe9),
	.dffe71(dffe7),
	.dffe81(dffe8),
	.dffe19(dffe1),
	.dffe21(dffe2),
	.dffe31(dffe3),
	.dffe41(dffe4),
	.dffe51(dffe5),
	.dffe61(dffe6),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module nco_test_add_sub_jdg_2 (
	a_17,
	xordvalue_12,
	a_16,
	a_15,
	a_14,
	a_13,
	a_12,
	a_11,
	xordvalue_11,
	a_10,
	xordvalue_10,
	a_9,
	xordvalue_9,
	a_8,
	xordvalue_8,
	a_7,
	xordvalue_7,
	a_6,
	xordvalue_6,
	a_5,
	xordvalue_5,
	a_0,
	xordvalue_0,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	a_4,
	xordvalue_4,
	dffe181,
	dffe171,
	dffe161,
	dffe151,
	dffe141,
	dffe131,
	dffe121,
	dffe111,
	dffe101,
	dffe91,
	dffe71,
	dffe81,
	dffe19,
	dffe21,
	dffe31,
	dffe41,
	dffe51,
	dffe61,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_12;
input 	a_16;
input 	a_15;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	xordvalue_11;
input 	a_10;
input 	xordvalue_10;
input 	a_9;
input 	xordvalue_9;
input 	a_8;
input 	xordvalue_8;
input 	a_7;
input 	xordvalue_7;
input 	a_6;
input 	xordvalue_6;
input 	a_5;
input 	xordvalue_5;
input 	a_0;
input 	xordvalue_0;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
input 	a_4;
input 	xordvalue_4;
output 	dffe181;
output 	dffe171;
output 	dffe161;
output 	dffe151;
output 	dffe141;
output 	dffe131;
output 	dffe121;
output 	dffe111;
output 	dffe101;
output 	dffe91;
output 	dffe71;
output 	dffe81;
output 	dffe19;
output 	dffe21;
output 	dffe31;
output 	dffe41;
output 	dffe51;
output 	dffe61;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~COUT ;
wire \add_sub_cella[12]~COUT ;
wire \add_sub_cella[13]~COUT ;
wire \add_sub_cella[14]~COUT ;
wire \add_sub_cella[15]~COUT ;
wire \add_sub_cella[16]~COUT ;
wire \add_sub_cella[17]~sumout ;
wire \add_sub_cella[16]~sumout ;
wire \add_sub_cella[15]~sumout ;
wire \add_sub_cella[14]~sumout ;
wire \add_sub_cella[13]~sumout ;
wire \add_sub_cella[12]~sumout ;
wire \add_sub_cella[11]~sumout ;
wire \add_sub_cella[10]~sumout ;
wire \add_sub_cella[9]~sumout ;
wire \add_sub_cella[8]~sumout ;
wire \add_sub_cella[6]~sumout ;
wire \add_sub_cella[7]~sumout ;
wire \add_sub_cella[0]~sumout ;
wire \add_sub_cella[1]~sumout ;
wire \add_sub_cella[2]~sumout ;
wire \add_sub_cella[3]~sumout ;
wire \add_sub_cella[4]~sumout ;
wire \add_sub_cella[5]~sumout ;


dffeas dffe18(
	.clk(clock),
	.d(\add_sub_cella[17]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe181),
	.prn(vcc));
defparam dffe18.is_wysiwyg = "true";
defparam dffe18.power_up = "low";

dffeas dffe17(
	.clk(clock),
	.d(\add_sub_cella[16]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe171),
	.prn(vcc));
defparam dffe17.is_wysiwyg = "true";
defparam dffe17.power_up = "low";

dffeas dffe16(
	.clk(clock),
	.d(\add_sub_cella[15]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe161),
	.prn(vcc));
defparam dffe16.is_wysiwyg = "true";
defparam dffe16.power_up = "low";

dffeas dffe15(
	.clk(clock),
	.d(\add_sub_cella[14]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe151),
	.prn(vcc));
defparam dffe15.is_wysiwyg = "true";
defparam dffe15.power_up = "low";

dffeas dffe14(
	.clk(clock),
	.d(\add_sub_cella[13]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe141),
	.prn(vcc));
defparam dffe14.is_wysiwyg = "true";
defparam dffe14.power_up = "low";

dffeas dffe13(
	.clk(clock),
	.d(\add_sub_cella[12]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe131),
	.prn(vcc));
defparam dffe13.is_wysiwyg = "true";
defparam dffe13.power_up = "low";

dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe19),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

arriav_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_1),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_2),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_3),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_4),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_5),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_6),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_7),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_8),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_9),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_11),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(\add_sub_cella[11]~COUT ),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[12] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_12),
	.datag(gnd),
	.cin(\add_sub_cella[11]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[12]~sumout ),
	.cout(\add_sub_cella[12]~COUT ),
	.shareout());
defparam \add_sub_cella[12] .extended_lut = "off";
defparam \add_sub_cella[12] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[12] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[13] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_12),
	.datag(gnd),
	.cin(\add_sub_cella[12]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[13]~sumout ),
	.cout(\add_sub_cella[13]~COUT ),
	.shareout());
defparam \add_sub_cella[13] .extended_lut = "off";
defparam \add_sub_cella[13] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[13] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[14] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_12),
	.datag(gnd),
	.cin(\add_sub_cella[13]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[14]~sumout ),
	.cout(\add_sub_cella[14]~COUT ),
	.shareout());
defparam \add_sub_cella[14] .extended_lut = "off";
defparam \add_sub_cella[14] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[14] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[15] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_12),
	.datag(gnd),
	.cin(\add_sub_cella[14]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[15]~sumout ),
	.cout(\add_sub_cella[15]~COUT ),
	.shareout());
defparam \add_sub_cella[15] .extended_lut = "off";
defparam \add_sub_cella[15] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[15] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[16] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_16),
	.datae(gnd),
	.dataf(!xordvalue_12),
	.datag(gnd),
	.cin(\add_sub_cella[15]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[16]~sumout ),
	.cout(\add_sub_cella[16]~COUT ),
	.shareout());
defparam \add_sub_cella[16] .extended_lut = "off";
defparam \add_sub_cella[16] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[16] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[17] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_17),
	.datae(gnd),
	.dataf(!xordvalue_12),
	.datag(gnd),
	.cin(\add_sub_cella[16]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[17]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[17] .extended_lut = "off";
defparam \add_sub_cella[17] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[17] .shared_arith = "off";

endmodule

module nco_test_cordic_sxor_1p_lpm_3 (
	sin_o_0,
	dffe18,
	dffe17,
	dffe16,
	pipeline_dffe_17,
	dffe161,
	dffe181,
	dffe15,
	dffe171,
	dffe14,
	pipeline_dffe_16,
	dffe162,
	dffe13,
	pipeline_dffe_15,
	dffe151,
	dffe12,
	pipeline_dffe_14,
	dffe141,
	dffe11,
	pipeline_dffe_13,
	dffe131,
	dffe10,
	pipeline_dffe_12,
	dffe8,
	dffe9,
	dffe121,
	pipeline_dffe_11,
	dffe111,
	dffe1,
	pipeline_dffe_10,
	dffe2,
	dffe3,
	dffe4,
	dffe5,
	dffe6,
	dffe7,
	dffe101,
	pipeline_dffe_9,
	dffe91,
	pipeline_dffe_8,
	dffe71,
	dffe81,
	pipeline_dffe_6,
	pipeline_dffe_7,
	dffe19,
	dffe21,
	dffe31,
	dffe41,
	dffe51,
	dffe61,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	sin_o_0;
output 	dffe18;
output 	dffe17;
input 	dffe16;
input 	pipeline_dffe_17;
output 	dffe161;
input 	dffe181;
output 	dffe15;
input 	dffe171;
output 	dffe14;
input 	pipeline_dffe_16;
input 	dffe162;
output 	dffe13;
input 	pipeline_dffe_15;
input 	dffe151;
output 	dffe12;
input 	pipeline_dffe_14;
input 	dffe141;
output 	dffe11;
input 	pipeline_dffe_13;
input 	dffe131;
output 	dffe10;
input 	pipeline_dffe_12;
output 	dffe8;
output 	dffe9;
input 	dffe121;
input 	pipeline_dffe_11;
input 	dffe111;
output 	dffe1;
input 	pipeline_dffe_10;
output 	dffe2;
output 	dffe3;
output 	dffe4;
output 	dffe5;
output 	dffe6;
output 	dffe7;
input 	dffe101;
input 	pipeline_dffe_9;
input 	dffe91;
input 	pipeline_dffe_8;
input 	dffe71;
input 	dffe81;
input 	pipeline_dffe_6;
input 	pipeline_dffe_7;
input 	dffe19;
input 	dffe21;
input 	dffe31;
input 	dffe41;
input 	dffe51;
input 	dffe61;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[17]~q ;
wire \xordvalue[11]~q ;
wire \Add0~1_sumout ;
wire \a[16]~q ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \a[15]~q ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \a[14]~q ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \a[13]~q ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \a[12]~q ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \a[11]~q ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \a[10]~q ;
wire \xordvalue[10]~q ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \a[9]~q ;
wire \xordvalue[9]~q ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \a[8]~q ;
wire \xordvalue[8]~q ;
wire \a[7]~q ;
wire \xordvalue[7]~q ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \a[6]~q ;
wire \xordvalue[6]~q ;
wire \a[0]~q ;
wire \xordvalue[0]~q ;
wire \a[1]~q ;
wire \xordvalue[1]~q ;
wire \a[2]~q ;
wire \xordvalue[2]~q ;
wire \a[3]~q ;
wire \xordvalue[3]~q ;
wire \a[4]~q ;
wire \xordvalue[4]~q ;
wire \a[5]~q ;
wire \xordvalue[5]~q ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~51 ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~55 ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~59 ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~63 ;
wire \Add0~65_sumout ;
wire \Add0~66 ;
wire \Add0~67 ;
wire \Add0~69_sumout ;
wire \Add0~70 ;
wire \Add0~71 ;
wire \xordvalue~0_combout ;
wire \xordvalue~1_combout ;
wire \xordvalue~2_combout ;
wire \xordvalue~3_combout ;
wire \xordvalue~4_combout ;
wire \xordvalue~5_combout ;
wire \xordvalue~6_combout ;
wire \xordvalue~7_combout ;
wire \xordvalue~8_combout ;
wire \xordvalue~9_combout ;
wire \xordvalue~10_combout ;
wire \xordvalue~11_combout ;


nco_test_lpm_add_sub_22 u0(
	.a_17(\a[17]~q ),
	.xordvalue_11(\xordvalue[11]~q ),
	.a_16(\a[16]~q ),
	.a_15(\a[15]~q ),
	.a_14(\a[14]~q ),
	.a_13(\a[13]~q ),
	.a_12(\a[12]~q ),
	.a_11(\a[11]~q ),
	.a_10(\a[10]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.a_9(\a[9]~q ),
	.xordvalue_9(\xordvalue[9]~q ),
	.a_8(\a[8]~q ),
	.xordvalue_8(\xordvalue[8]~q ),
	.a_7(\a[7]~q ),
	.xordvalue_7(\xordvalue[7]~q ),
	.a_6(\a[6]~q ),
	.xordvalue_6(\xordvalue[6]~q ),
	.a_0(\a[0]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_1(\a[1]~q ),
	.xordvalue_1(\xordvalue[1]~q ),
	.a_2(\a[2]~q ),
	.xordvalue_2(\xordvalue[2]~q ),
	.a_3(\a[3]~q ),
	.xordvalue_3(\xordvalue[3]~q ),
	.a_4(\a[4]~q ),
	.xordvalue_4(\xordvalue[4]~q ),
	.a_5(\a[5]~q ),
	.xordvalue_5(\xordvalue[5]~q ),
	.dffe18(dffe18),
	.dffe17(dffe17),
	.dffe16(dffe161),
	.dffe15(dffe15),
	.dffe14(dffe14),
	.dffe13(dffe13),
	.dffe12(dffe12),
	.dffe11(dffe11),
	.dffe10(dffe10),
	.dffe8(dffe8),
	.dffe9(dffe9),
	.dffe1(dffe1),
	.dffe2(dffe2),
	.dffe3(dffe3),
	.dffe4(dffe4),
	.dffe5(dffe5),
	.dffe6(dffe6),
	.dffe7(dffe7),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[17] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[17]~q ),
	.prn(vcc));
defparam \a[17] .is_wysiwyg = "true";
defparam \a[17] .power_up = "low";

dffeas \xordvalue[11] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[11]~q ),
	.prn(vcc));
defparam \xordvalue[11] .is_wysiwyg = "true";
defparam \xordvalue[11] .power_up = "low";

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe181),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "on";

dffeas \a[16] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[16]~q ),
	.prn(vcc));
defparam \a[16] .is_wysiwyg = "true";
defparam \a[16] .power_up = "low";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe171),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~5 .shared_arith = "on";

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe162),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~9 .shared_arith = "on";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~13 .shared_arith = "on";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~17 .shared_arith = "on";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "on";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~25 .shared_arith = "on";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(\xordvalue~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~29 .shared_arith = "on";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \xordvalue[9] (
	.clk(clk),
	.d(\xordvalue~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[9]~q ),
	.prn(vcc));
defparam \xordvalue[9] .is_wysiwyg = "true";
defparam \xordvalue[9] .power_up = "low";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~33 .shared_arith = "on";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \xordvalue[8] (
	.clk(clk),
	.d(\xordvalue~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[8]~q ),
	.prn(vcc));
defparam \xordvalue[8] .is_wysiwyg = "true";
defparam \xordvalue[8] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \xordvalue[7] (
	.clk(clk),
	.d(\xordvalue~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[7]~q ),
	.prn(vcc));
defparam \xordvalue[7] .is_wysiwyg = "true";
defparam \xordvalue[7] .power_up = "low";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~37 .shared_arith = "on";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(\Add0~47 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~41 .shared_arith = "on";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \xordvalue[6] (
	.clk(clk),
	.d(\xordvalue~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[6]~q ),
	.prn(vcc));
defparam \xordvalue[6] .is_wysiwyg = "true";
defparam \xordvalue[6] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \xordvalue[1] (
	.clk(clk),
	.d(\xordvalue~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[1]~q ),
	.prn(vcc));
defparam \xordvalue[1] .is_wysiwyg = "true";
defparam \xordvalue[1] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \xordvalue[2] (
	.clk(clk),
	.d(\xordvalue~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[2]~q ),
	.prn(vcc));
defparam \xordvalue[2] .is_wysiwyg = "true";
defparam \xordvalue[2] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \xordvalue[3] (
	.clk(clk),
	.d(\xordvalue~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[3]~q ),
	.prn(vcc));
defparam \xordvalue[3] .is_wysiwyg = "true";
defparam \xordvalue[3] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \xordvalue[4] (
	.clk(clk),
	.d(\xordvalue~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[4]~q ),
	.prn(vcc));
defparam \xordvalue[4] .is_wysiwyg = "true";
defparam \xordvalue[4] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \xordvalue[5] (
	.clk(clk),
	.d(\xordvalue~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[5]~q ),
	.prn(vcc));
defparam \xordvalue[5] .is_wysiwyg = "true";
defparam \xordvalue[5] .power_up = "low";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~70 ),
	.sharein(\Add0~71 ),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout(\Add0~47 ));
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~45 .shared_arith = "on";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!dffe19),
	.datad(!dffe16),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout(\Add0~51 ));
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add0~49 .shared_arith = "on";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(\Add0~51 ),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout(\Add0~55 ));
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~53 .shared_arith = "on";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(\Add0~55 ),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout(\Add0~59 ));
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~57 .shared_arith = "on";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(\Add0~59 ),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout(\Add0~63 ));
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~61 .shared_arith = "on";

arriav_lcell_comb \Add0~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(\Add0~63 ),
	.combout(),
	.sumout(\Add0~65_sumout ),
	.cout(\Add0~66 ),
	.shareout(\Add0~67 ));
defparam \Add0~65 .extended_lut = "off";
defparam \Add0~65 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~65 .shared_arith = "on";

arriav_lcell_comb \Add0~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~66 ),
	.sharein(\Add0~67 ),
	.combout(),
	.sumout(\Add0~69_sumout ),
	.cout(\Add0~70 ),
	.shareout(\Add0~71 ));
defparam \Add0~69 .extended_lut = "off";
defparam \Add0~69 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~69 .shared_arith = "on";

arriav_lcell_comb \xordvalue~0 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_17),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

arriav_lcell_comb \xordvalue~1 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~1 .extended_lut = "off";
defparam \xordvalue~1 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~1 .shared_arith = "off";

arriav_lcell_comb \xordvalue~2 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_15),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~2 .extended_lut = "off";
defparam \xordvalue~2 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~2 .shared_arith = "off";

arriav_lcell_comb \xordvalue~3 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_14),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~3 .extended_lut = "off";
defparam \xordvalue~3 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~3 .shared_arith = "off";

arriav_lcell_comb \xordvalue~4 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_13),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~4 .extended_lut = "off";
defparam \xordvalue~4 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~4 .shared_arith = "off";

arriav_lcell_comb \xordvalue~5 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_12),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~5 .extended_lut = "off";
defparam \xordvalue~5 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~5 .shared_arith = "off";

arriav_lcell_comb \xordvalue~6 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_6),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~6 .extended_lut = "off";
defparam \xordvalue~6 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~6 .shared_arith = "off";

arriav_lcell_comb \xordvalue~7 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_7),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~7 .extended_lut = "off";
defparam \xordvalue~7 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~7 .shared_arith = "off";

arriav_lcell_comb \xordvalue~8 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_8),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~8 .extended_lut = "off";
defparam \xordvalue~8 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~8 .shared_arith = "off";

arriav_lcell_comb \xordvalue~9 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_9),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~9 .extended_lut = "off";
defparam \xordvalue~9 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~9 .shared_arith = "off";

arriav_lcell_comb \xordvalue~10 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_10),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~10 .extended_lut = "off";
defparam \xordvalue~10 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~10 .shared_arith = "off";

arriav_lcell_comb \xordvalue~11 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_11),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~11 .extended_lut = "off";
defparam \xordvalue~11 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~11 .shared_arith = "off";

endmodule

module nco_test_lpm_add_sub_22 (
	a_17,
	xordvalue_11,
	a_16,
	a_15,
	a_14,
	a_13,
	a_12,
	a_11,
	a_10,
	xordvalue_10,
	a_9,
	xordvalue_9,
	a_8,
	xordvalue_8,
	a_7,
	xordvalue_7,
	a_6,
	xordvalue_6,
	a_0,
	xordvalue_0,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	a_4,
	xordvalue_4,
	a_5,
	xordvalue_5,
	dffe18,
	dffe17,
	dffe16,
	dffe15,
	dffe14,
	dffe13,
	dffe12,
	dffe11,
	dffe10,
	dffe8,
	dffe9,
	dffe1,
	dffe2,
	dffe3,
	dffe4,
	dffe5,
	dffe6,
	dffe7,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_11;
input 	a_16;
input 	a_15;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_10;
input 	xordvalue_10;
input 	a_9;
input 	xordvalue_9;
input 	a_8;
input 	xordvalue_8;
input 	a_7;
input 	xordvalue_7;
input 	a_6;
input 	xordvalue_6;
input 	a_0;
input 	xordvalue_0;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
input 	a_4;
input 	xordvalue_4;
input 	a_5;
input 	xordvalue_5;
output 	dffe18;
output 	dffe17;
output 	dffe16;
output 	dffe15;
output 	dffe14;
output 	dffe13;
output 	dffe12;
output 	dffe11;
output 	dffe10;
output 	dffe8;
output 	dffe9;
output 	dffe1;
output 	dffe2;
output 	dffe3;
output 	dffe4;
output 	dffe5;
output 	dffe6;
output 	dffe7;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_add_sub_jdg_3 auto_generated(
	.a_17(a_17),
	.xordvalue_11(xordvalue_11),
	.a_16(a_16),
	.a_15(a_15),
	.a_14(a_14),
	.a_13(a_13),
	.a_12(a_12),
	.a_11(a_11),
	.a_10(a_10),
	.xordvalue_10(xordvalue_10),
	.a_9(a_9),
	.xordvalue_9(xordvalue_9),
	.a_8(a_8),
	.xordvalue_8(xordvalue_8),
	.a_7(a_7),
	.xordvalue_7(xordvalue_7),
	.a_6(a_6),
	.xordvalue_6(xordvalue_6),
	.a_0(a_0),
	.xordvalue_0(xordvalue_0),
	.a_1(a_1),
	.xordvalue_1(xordvalue_1),
	.a_2(a_2),
	.xordvalue_2(xordvalue_2),
	.a_3(a_3),
	.xordvalue_3(xordvalue_3),
	.a_4(a_4),
	.xordvalue_4(xordvalue_4),
	.a_5(a_5),
	.xordvalue_5(xordvalue_5),
	.dffe181(dffe18),
	.dffe171(dffe17),
	.dffe161(dffe16),
	.dffe151(dffe15),
	.dffe141(dffe14),
	.dffe131(dffe13),
	.dffe121(dffe12),
	.dffe111(dffe11),
	.dffe101(dffe10),
	.dffe81(dffe8),
	.dffe91(dffe9),
	.dffe19(dffe1),
	.dffe21(dffe2),
	.dffe31(dffe3),
	.dffe41(dffe4),
	.dffe51(dffe5),
	.dffe61(dffe6),
	.dffe71(dffe7),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module nco_test_add_sub_jdg_3 (
	a_17,
	xordvalue_11,
	a_16,
	a_15,
	a_14,
	a_13,
	a_12,
	a_11,
	a_10,
	xordvalue_10,
	a_9,
	xordvalue_9,
	a_8,
	xordvalue_8,
	a_7,
	xordvalue_7,
	a_6,
	xordvalue_6,
	a_0,
	xordvalue_0,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	a_4,
	xordvalue_4,
	a_5,
	xordvalue_5,
	dffe181,
	dffe171,
	dffe161,
	dffe151,
	dffe141,
	dffe131,
	dffe121,
	dffe111,
	dffe101,
	dffe81,
	dffe91,
	dffe19,
	dffe21,
	dffe31,
	dffe41,
	dffe51,
	dffe61,
	dffe71,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_11;
input 	a_16;
input 	a_15;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_10;
input 	xordvalue_10;
input 	a_9;
input 	xordvalue_9;
input 	a_8;
input 	xordvalue_8;
input 	a_7;
input 	xordvalue_7;
input 	a_6;
input 	xordvalue_6;
input 	a_0;
input 	xordvalue_0;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
input 	a_4;
input 	xordvalue_4;
input 	a_5;
input 	xordvalue_5;
output 	dffe181;
output 	dffe171;
output 	dffe161;
output 	dffe151;
output 	dffe141;
output 	dffe131;
output 	dffe121;
output 	dffe111;
output 	dffe101;
output 	dffe81;
output 	dffe91;
output 	dffe19;
output 	dffe21;
output 	dffe31;
output 	dffe41;
output 	dffe51;
output 	dffe61;
output 	dffe71;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~COUT ;
wire \add_sub_cella[12]~COUT ;
wire \add_sub_cella[13]~COUT ;
wire \add_sub_cella[14]~COUT ;
wire \add_sub_cella[15]~COUT ;
wire \add_sub_cella[16]~COUT ;
wire \add_sub_cella[17]~sumout ;
wire \add_sub_cella[16]~sumout ;
wire \add_sub_cella[15]~sumout ;
wire \add_sub_cella[14]~sumout ;
wire \add_sub_cella[13]~sumout ;
wire \add_sub_cella[12]~sumout ;
wire \add_sub_cella[11]~sumout ;
wire \add_sub_cella[10]~sumout ;
wire \add_sub_cella[9]~sumout ;
wire \add_sub_cella[7]~sumout ;
wire \add_sub_cella[8]~sumout ;
wire \add_sub_cella[0]~sumout ;
wire \add_sub_cella[1]~sumout ;
wire \add_sub_cella[2]~sumout ;
wire \add_sub_cella[3]~sumout ;
wire \add_sub_cella[4]~sumout ;
wire \add_sub_cella[5]~sumout ;
wire \add_sub_cella[6]~sumout ;


dffeas dffe18(
	.clk(clock),
	.d(\add_sub_cella[17]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe181),
	.prn(vcc));
defparam dffe18.is_wysiwyg = "true";
defparam dffe18.power_up = "low";

dffeas dffe17(
	.clk(clock),
	.d(\add_sub_cella[16]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe171),
	.prn(vcc));
defparam dffe17.is_wysiwyg = "true";
defparam dffe17.power_up = "low";

dffeas dffe16(
	.clk(clock),
	.d(\add_sub_cella[15]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe161),
	.prn(vcc));
defparam dffe16.is_wysiwyg = "true";
defparam dffe16.power_up = "low";

dffeas dffe15(
	.clk(clock),
	.d(\add_sub_cella[14]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe151),
	.prn(vcc));
defparam dffe15.is_wysiwyg = "true";
defparam dffe15.power_up = "low";

dffeas dffe14(
	.clk(clock),
	.d(\add_sub_cella[13]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe141),
	.prn(vcc));
defparam dffe14.is_wysiwyg = "true";
defparam dffe14.power_up = "low";

dffeas dffe13(
	.clk(clock),
	.d(\add_sub_cella[12]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe131),
	.prn(vcc));
defparam dffe13.is_wysiwyg = "true";
defparam dffe13.power_up = "low";

dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe19),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

arriav_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_1),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_2),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_3),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_4),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_5),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_6),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_7),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_8),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_9),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_11),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(\add_sub_cella[11]~COUT ),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[12] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_11),
	.datag(gnd),
	.cin(\add_sub_cella[11]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[12]~sumout ),
	.cout(\add_sub_cella[12]~COUT ),
	.shareout());
defparam \add_sub_cella[12] .extended_lut = "off";
defparam \add_sub_cella[12] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[12] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[13] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_11),
	.datag(gnd),
	.cin(\add_sub_cella[12]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[13]~sumout ),
	.cout(\add_sub_cella[13]~COUT ),
	.shareout());
defparam \add_sub_cella[13] .extended_lut = "off";
defparam \add_sub_cella[13] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[13] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[14] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_11),
	.datag(gnd),
	.cin(\add_sub_cella[13]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[14]~sumout ),
	.cout(\add_sub_cella[14]~COUT ),
	.shareout());
defparam \add_sub_cella[14] .extended_lut = "off";
defparam \add_sub_cella[14] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[14] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[15] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_11),
	.datag(gnd),
	.cin(\add_sub_cella[14]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[15]~sumout ),
	.cout(\add_sub_cella[15]~COUT ),
	.shareout());
defparam \add_sub_cella[15] .extended_lut = "off";
defparam \add_sub_cella[15] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[15] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[16] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_16),
	.datae(gnd),
	.dataf(!xordvalue_11),
	.datag(gnd),
	.cin(\add_sub_cella[15]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[16]~sumout ),
	.cout(\add_sub_cella[16]~COUT ),
	.shareout());
defparam \add_sub_cella[16] .extended_lut = "off";
defparam \add_sub_cella[16] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[16] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[17] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_17),
	.datae(gnd),
	.dataf(!xordvalue_11),
	.datag(gnd),
	.cin(\add_sub_cella[16]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[17]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[17] .extended_lut = "off";
defparam \add_sub_cella[17] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[17] .shared_arith = "off";

endmodule

module nco_test_cordic_sxor_1p_lpm_4 (
	sin_o_0,
	dffe18,
	dffe17,
	dffe16,
	dffe161,
	dffe181,
	pipeline_dffe_17,
	dffe15,
	dffe14,
	pipeline_dffe_16,
	dffe171,
	dffe13,
	pipeline_dffe_15,
	dffe162,
	dffe12,
	pipeline_dffe_14,
	dffe151,
	dffe11,
	pipeline_dffe_13,
	dffe141,
	dffe9,
	dffe10,
	pipeline_dffe_12,
	dffe131,
	pipeline_dffe_11,
	dffe1,
	dffe121,
	dffe2,
	dffe3,
	dffe4,
	dffe5,
	dffe6,
	dffe7,
	dffe8,
	pipeline_dffe_10,
	dffe111,
	pipeline_dffe_9,
	dffe101,
	dffe81,
	dffe91,
	pipeline_dffe_8,
	pipeline_dffe_7,
	dffe19,
	dffe21,
	dffe31,
	dffe41,
	dffe51,
	dffe61,
	dffe71,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	sin_o_0;
output 	dffe18;
output 	dffe17;
input 	dffe16;
output 	dffe161;
input 	dffe181;
input 	pipeline_dffe_17;
output 	dffe15;
output 	dffe14;
input 	pipeline_dffe_16;
input 	dffe171;
output 	dffe13;
input 	pipeline_dffe_15;
input 	dffe162;
output 	dffe12;
input 	pipeline_dffe_14;
input 	dffe151;
output 	dffe11;
input 	pipeline_dffe_13;
input 	dffe141;
output 	dffe9;
output 	dffe10;
input 	pipeline_dffe_12;
input 	dffe131;
input 	pipeline_dffe_11;
output 	dffe1;
input 	dffe121;
output 	dffe2;
output 	dffe3;
output 	dffe4;
output 	dffe5;
output 	dffe6;
output 	dffe7;
output 	dffe8;
input 	pipeline_dffe_10;
input 	dffe111;
input 	pipeline_dffe_9;
input 	dffe101;
input 	dffe81;
input 	dffe91;
input 	pipeline_dffe_8;
input 	pipeline_dffe_7;
input 	dffe19;
input 	dffe21;
input 	dffe31;
input 	dffe41;
input 	dffe51;
input 	dffe61;
input 	dffe71;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[17]~q ;
wire \xordvalue[10]~q ;
wire \Add0~1_sumout ;
wire \a[16]~q ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \a[15]~q ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \a[14]~q ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \a[13]~q ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \a[12]~q ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \a[11]~q ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \a[10]~q ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \a[9]~q ;
wire \xordvalue[9]~q ;
wire \a[8]~q ;
wire \xordvalue[8]~q ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \a[7]~q ;
wire \xordvalue[7]~q ;
wire \a[0]~q ;
wire \xordvalue[0]~q ;
wire \a[1]~q ;
wire \xordvalue[1]~q ;
wire \a[2]~q ;
wire \xordvalue[2]~q ;
wire \a[3]~q ;
wire \xordvalue[3]~q ;
wire \a[4]~q ;
wire \xordvalue[4]~q ;
wire \a[5]~q ;
wire \xordvalue[5]~q ;
wire \a[6]~q ;
wire \xordvalue[6]~q ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~51 ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~55 ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~59 ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~63 ;
wire \Add0~65_sumout ;
wire \Add0~66 ;
wire \Add0~67 ;
wire \Add0~69_sumout ;
wire \Add0~70 ;
wire \Add0~71 ;
wire \xordvalue~0_combout ;
wire \xordvalue~1_combout ;
wire \xordvalue~2_combout ;
wire \xordvalue~3_combout ;
wire \xordvalue~4_combout ;
wire \xordvalue~5_combout ;
wire \xordvalue~6_combout ;
wire \xordvalue~7_combout ;
wire \xordvalue~8_combout ;
wire \xordvalue~9_combout ;
wire \xordvalue~10_combout ;


nco_test_lpm_add_sub_23 u0(
	.a_17(\a[17]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.a_16(\a[16]~q ),
	.a_15(\a[15]~q ),
	.a_14(\a[14]~q ),
	.a_13(\a[13]~q ),
	.a_12(\a[12]~q ),
	.a_11(\a[11]~q ),
	.a_10(\a[10]~q ),
	.a_9(\a[9]~q ),
	.xordvalue_9(\xordvalue[9]~q ),
	.a_8(\a[8]~q ),
	.xordvalue_8(\xordvalue[8]~q ),
	.a_7(\a[7]~q ),
	.xordvalue_7(\xordvalue[7]~q ),
	.a_0(\a[0]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_1(\a[1]~q ),
	.xordvalue_1(\xordvalue[1]~q ),
	.a_2(\a[2]~q ),
	.xordvalue_2(\xordvalue[2]~q ),
	.a_3(\a[3]~q ),
	.xordvalue_3(\xordvalue[3]~q ),
	.a_4(\a[4]~q ),
	.xordvalue_4(\xordvalue[4]~q ),
	.a_5(\a[5]~q ),
	.xordvalue_5(\xordvalue[5]~q ),
	.a_6(\a[6]~q ),
	.xordvalue_6(\xordvalue[6]~q ),
	.dffe18(dffe18),
	.dffe17(dffe17),
	.dffe16(dffe161),
	.dffe15(dffe15),
	.dffe14(dffe14),
	.dffe13(dffe13),
	.dffe12(dffe12),
	.dffe11(dffe11),
	.dffe9(dffe9),
	.dffe10(dffe10),
	.dffe1(dffe1),
	.dffe2(dffe2),
	.dffe3(dffe3),
	.dffe4(dffe4),
	.dffe5(dffe5),
	.dffe6(dffe6),
	.dffe7(dffe7),
	.dffe8(dffe8),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[17] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[17]~q ),
	.prn(vcc));
defparam \a[17] .is_wysiwyg = "true";
defparam \a[17] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe181),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "on";

dffeas \a[16] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[16]~q ),
	.prn(vcc));
defparam \a[16] .is_wysiwyg = "true";
defparam \a[16] .power_up = "low";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe171),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~5 .shared_arith = "on";

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe162),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~9 .shared_arith = "on";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~13 .shared_arith = "on";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~17 .shared_arith = "on";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "on";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~25 .shared_arith = "on";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~29 .shared_arith = "on";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \xordvalue[9] (
	.clk(clk),
	.d(\xordvalue~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[9]~q ),
	.prn(vcc));
defparam \xordvalue[9] .is_wysiwyg = "true";
defparam \xordvalue[9] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \xordvalue[8] (
	.clk(clk),
	.d(\xordvalue~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[8]~q ),
	.prn(vcc));
defparam \xordvalue[8] .is_wysiwyg = "true";
defparam \xordvalue[8] .power_up = "low";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~33 .shared_arith = "on";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~37 .shared_arith = "on";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \xordvalue[7] (
	.clk(clk),
	.d(\xordvalue~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[7]~q ),
	.prn(vcc));
defparam \xordvalue[7] .is_wysiwyg = "true";
defparam \xordvalue[7] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \xordvalue[1] (
	.clk(clk),
	.d(\xordvalue~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[1]~q ),
	.prn(vcc));
defparam \xordvalue[1] .is_wysiwyg = "true";
defparam \xordvalue[1] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \xordvalue[2] (
	.clk(clk),
	.d(\xordvalue~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[2]~q ),
	.prn(vcc));
defparam \xordvalue[2] .is_wysiwyg = "true";
defparam \xordvalue[2] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \xordvalue[3] (
	.clk(clk),
	.d(\xordvalue~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[3]~q ),
	.prn(vcc));
defparam \xordvalue[3] .is_wysiwyg = "true";
defparam \xordvalue[3] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \xordvalue[4] (
	.clk(clk),
	.d(\xordvalue~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[4]~q ),
	.prn(vcc));
defparam \xordvalue[4] .is_wysiwyg = "true";
defparam \xordvalue[4] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \xordvalue[5] (
	.clk(clk),
	.d(\xordvalue~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[5]~q ),
	.prn(vcc));
defparam \xordvalue[5] .is_wysiwyg = "true";
defparam \xordvalue[5] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \xordvalue[6] (
	.clk(clk),
	.d(\xordvalue~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[6]~q ),
	.prn(vcc));
defparam \xordvalue[6] .is_wysiwyg = "true";
defparam \xordvalue[6] .power_up = "low";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~70 ),
	.sharein(\Add0~71 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~41 .shared_arith = "on";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!dffe19),
	.datad(!dffe16),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout(\Add0~47 ));
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add0~45 .shared_arith = "on";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(\Add0~47 ),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout(\Add0~51 ));
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~49 .shared_arith = "on";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(\Add0~51 ),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout(\Add0~55 ));
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~53 .shared_arith = "on";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(\Add0~55 ),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout(\Add0~59 ));
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~57 .shared_arith = "on";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(\Add0~59 ),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout(\Add0~63 ));
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~61 .shared_arith = "on";

arriav_lcell_comb \Add0~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(\Add0~63 ),
	.combout(),
	.sumout(\Add0~65_sumout ),
	.cout(\Add0~66 ),
	.shareout(\Add0~67 ));
defparam \Add0~65 .extended_lut = "off";
defparam \Add0~65 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~65 .shared_arith = "on";

arriav_lcell_comb \Add0~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~66 ),
	.sharein(\Add0~67 ),
	.combout(),
	.sumout(\Add0~69_sumout ),
	.cout(\Add0~70 ),
	.shareout(\Add0~71 ));
defparam \Add0~69 .extended_lut = "off";
defparam \Add0~69 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~69 .shared_arith = "on";

arriav_lcell_comb \xordvalue~0 (
	.dataa(!pipeline_dffe_17),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

arriav_lcell_comb \xordvalue~1 (
	.dataa(!pipeline_dffe_16),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~1 .extended_lut = "off";
defparam \xordvalue~1 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~1 .shared_arith = "off";

arriav_lcell_comb \xordvalue~2 (
	.dataa(!pipeline_dffe_15),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~2 .extended_lut = "off";
defparam \xordvalue~2 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~2 .shared_arith = "off";

arriav_lcell_comb \xordvalue~3 (
	.dataa(!pipeline_dffe_14),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~3 .extended_lut = "off";
defparam \xordvalue~3 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~3 .shared_arith = "off";

arriav_lcell_comb \xordvalue~4 (
	.dataa(!pipeline_dffe_7),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~4 .extended_lut = "off";
defparam \xordvalue~4 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~4 .shared_arith = "off";

arriav_lcell_comb \xordvalue~5 (
	.dataa(!pipeline_dffe_8),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~5 .extended_lut = "off";
defparam \xordvalue~5 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~5 .shared_arith = "off";

arriav_lcell_comb \xordvalue~6 (
	.dataa(!pipeline_dffe_9),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~6 .extended_lut = "off";
defparam \xordvalue~6 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~6 .shared_arith = "off";

arriav_lcell_comb \xordvalue~7 (
	.dataa(!pipeline_dffe_10),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~7 .extended_lut = "off";
defparam \xordvalue~7 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~7 .shared_arith = "off";

arriav_lcell_comb \xordvalue~8 (
	.dataa(!pipeline_dffe_11),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~8 .extended_lut = "off";
defparam \xordvalue~8 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~8 .shared_arith = "off";

arriav_lcell_comb \xordvalue~9 (
	.dataa(!pipeline_dffe_12),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~9 .extended_lut = "off";
defparam \xordvalue~9 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~9 .shared_arith = "off";

arriav_lcell_comb \xordvalue~10 (
	.dataa(!pipeline_dffe_13),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~10 .extended_lut = "off";
defparam \xordvalue~10 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~10 .shared_arith = "off";

endmodule

module nco_test_lpm_add_sub_23 (
	a_17,
	xordvalue_10,
	a_16,
	a_15,
	a_14,
	a_13,
	a_12,
	a_11,
	a_10,
	a_9,
	xordvalue_9,
	a_8,
	xordvalue_8,
	a_7,
	xordvalue_7,
	a_0,
	xordvalue_0,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	a_4,
	xordvalue_4,
	a_5,
	xordvalue_5,
	a_6,
	xordvalue_6,
	dffe18,
	dffe17,
	dffe16,
	dffe15,
	dffe14,
	dffe13,
	dffe12,
	dffe11,
	dffe9,
	dffe10,
	dffe1,
	dffe2,
	dffe3,
	dffe4,
	dffe5,
	dffe6,
	dffe7,
	dffe8,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_10;
input 	a_16;
input 	a_15;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_10;
input 	a_9;
input 	xordvalue_9;
input 	a_8;
input 	xordvalue_8;
input 	a_7;
input 	xordvalue_7;
input 	a_0;
input 	xordvalue_0;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
input 	a_4;
input 	xordvalue_4;
input 	a_5;
input 	xordvalue_5;
input 	a_6;
input 	xordvalue_6;
output 	dffe18;
output 	dffe17;
output 	dffe16;
output 	dffe15;
output 	dffe14;
output 	dffe13;
output 	dffe12;
output 	dffe11;
output 	dffe9;
output 	dffe10;
output 	dffe1;
output 	dffe2;
output 	dffe3;
output 	dffe4;
output 	dffe5;
output 	dffe6;
output 	dffe7;
output 	dffe8;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_add_sub_jdg_4 auto_generated(
	.a_17(a_17),
	.xordvalue_10(xordvalue_10),
	.a_16(a_16),
	.a_15(a_15),
	.a_14(a_14),
	.a_13(a_13),
	.a_12(a_12),
	.a_11(a_11),
	.a_10(a_10),
	.a_9(a_9),
	.xordvalue_9(xordvalue_9),
	.a_8(a_8),
	.xordvalue_8(xordvalue_8),
	.a_7(a_7),
	.xordvalue_7(xordvalue_7),
	.a_0(a_0),
	.xordvalue_0(xordvalue_0),
	.a_1(a_1),
	.xordvalue_1(xordvalue_1),
	.a_2(a_2),
	.xordvalue_2(xordvalue_2),
	.a_3(a_3),
	.xordvalue_3(xordvalue_3),
	.a_4(a_4),
	.xordvalue_4(xordvalue_4),
	.a_5(a_5),
	.xordvalue_5(xordvalue_5),
	.a_6(a_6),
	.xordvalue_6(xordvalue_6),
	.dffe181(dffe18),
	.dffe171(dffe17),
	.dffe161(dffe16),
	.dffe151(dffe15),
	.dffe141(dffe14),
	.dffe131(dffe13),
	.dffe121(dffe12),
	.dffe111(dffe11),
	.dffe91(dffe9),
	.dffe101(dffe10),
	.dffe19(dffe1),
	.dffe21(dffe2),
	.dffe31(dffe3),
	.dffe41(dffe4),
	.dffe51(dffe5),
	.dffe61(dffe6),
	.dffe71(dffe7),
	.dffe81(dffe8),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module nco_test_add_sub_jdg_4 (
	a_17,
	xordvalue_10,
	a_16,
	a_15,
	a_14,
	a_13,
	a_12,
	a_11,
	a_10,
	a_9,
	xordvalue_9,
	a_8,
	xordvalue_8,
	a_7,
	xordvalue_7,
	a_0,
	xordvalue_0,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	a_4,
	xordvalue_4,
	a_5,
	xordvalue_5,
	a_6,
	xordvalue_6,
	dffe181,
	dffe171,
	dffe161,
	dffe151,
	dffe141,
	dffe131,
	dffe121,
	dffe111,
	dffe91,
	dffe101,
	dffe19,
	dffe21,
	dffe31,
	dffe41,
	dffe51,
	dffe61,
	dffe71,
	dffe81,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_10;
input 	a_16;
input 	a_15;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_10;
input 	a_9;
input 	xordvalue_9;
input 	a_8;
input 	xordvalue_8;
input 	a_7;
input 	xordvalue_7;
input 	a_0;
input 	xordvalue_0;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
input 	a_4;
input 	xordvalue_4;
input 	a_5;
input 	xordvalue_5;
input 	a_6;
input 	xordvalue_6;
output 	dffe181;
output 	dffe171;
output 	dffe161;
output 	dffe151;
output 	dffe141;
output 	dffe131;
output 	dffe121;
output 	dffe111;
output 	dffe91;
output 	dffe101;
output 	dffe19;
output 	dffe21;
output 	dffe31;
output 	dffe41;
output 	dffe51;
output 	dffe61;
output 	dffe71;
output 	dffe81;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~COUT ;
wire \add_sub_cella[12]~COUT ;
wire \add_sub_cella[13]~COUT ;
wire \add_sub_cella[14]~COUT ;
wire \add_sub_cella[15]~COUT ;
wire \add_sub_cella[16]~COUT ;
wire \add_sub_cella[17]~sumout ;
wire \add_sub_cella[16]~sumout ;
wire \add_sub_cella[15]~sumout ;
wire \add_sub_cella[14]~sumout ;
wire \add_sub_cella[13]~sumout ;
wire \add_sub_cella[12]~sumout ;
wire \add_sub_cella[11]~sumout ;
wire \add_sub_cella[10]~sumout ;
wire \add_sub_cella[8]~sumout ;
wire \add_sub_cella[9]~sumout ;
wire \add_sub_cella[0]~sumout ;
wire \add_sub_cella[1]~sumout ;
wire \add_sub_cella[2]~sumout ;
wire \add_sub_cella[3]~sumout ;
wire \add_sub_cella[4]~sumout ;
wire \add_sub_cella[5]~sumout ;
wire \add_sub_cella[6]~sumout ;
wire \add_sub_cella[7]~sumout ;


dffeas dffe18(
	.clk(clock),
	.d(\add_sub_cella[17]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe181),
	.prn(vcc));
defparam dffe18.is_wysiwyg = "true";
defparam dffe18.power_up = "low";

dffeas dffe17(
	.clk(clock),
	.d(\add_sub_cella[16]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe171),
	.prn(vcc));
defparam dffe17.is_wysiwyg = "true";
defparam dffe17.power_up = "low";

dffeas dffe16(
	.clk(clock),
	.d(\add_sub_cella[15]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe161),
	.prn(vcc));
defparam dffe16.is_wysiwyg = "true";
defparam dffe16.power_up = "low";

dffeas dffe15(
	.clk(clock),
	.d(\add_sub_cella[14]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe151),
	.prn(vcc));
defparam dffe15.is_wysiwyg = "true";
defparam dffe15.power_up = "low";

dffeas dffe14(
	.clk(clock),
	.d(\add_sub_cella[13]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe141),
	.prn(vcc));
defparam dffe14.is_wysiwyg = "true";
defparam dffe14.power_up = "low";

dffeas dffe13(
	.clk(clock),
	.d(\add_sub_cella[12]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe131),
	.prn(vcc));
defparam dffe13.is_wysiwyg = "true";
defparam dffe13.power_up = "low";

dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe19),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

arriav_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_1),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_2),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_3),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_4),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_5),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_6),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_7),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_8),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_9),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(\add_sub_cella[11]~COUT ),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[12] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[11]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[12]~sumout ),
	.cout(\add_sub_cella[12]~COUT ),
	.shareout());
defparam \add_sub_cella[12] .extended_lut = "off";
defparam \add_sub_cella[12] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[12] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[13] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[12]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[13]~sumout ),
	.cout(\add_sub_cella[13]~COUT ),
	.shareout());
defparam \add_sub_cella[13] .extended_lut = "off";
defparam \add_sub_cella[13] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[13] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[14] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[13]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[14]~sumout ),
	.cout(\add_sub_cella[14]~COUT ),
	.shareout());
defparam \add_sub_cella[14] .extended_lut = "off";
defparam \add_sub_cella[14] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[14] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[15] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[14]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[15]~sumout ),
	.cout(\add_sub_cella[15]~COUT ),
	.shareout());
defparam \add_sub_cella[15] .extended_lut = "off";
defparam \add_sub_cella[15] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[15] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[16] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_16),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[15]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[16]~sumout ),
	.cout(\add_sub_cella[16]~COUT ),
	.shareout());
defparam \add_sub_cella[16] .extended_lut = "off";
defparam \add_sub_cella[16] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[16] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[17] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_17),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[16]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[17]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[17] .extended_lut = "off";
defparam \add_sub_cella[17] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[17] .shared_arith = "off";

endmodule

module nco_test_cordic_sxor_1p_lpm_5 (
	sin_o_0,
	dffe18,
	dffe17,
	dffe16,
	pipeline_dffe_17,
	dffe161,
	dffe181,
	dffe15,
	dffe171,
	dffe14,
	pipeline_dffe_16,
	dffe162,
	dffe13,
	pipeline_dffe_15,
	dffe151,
	dffe12,
	pipeline_dffe_14,
	dffe10,
	dffe11,
	dffe141,
	pipeline_dffe_13,
	dffe131,
	dffe1,
	pipeline_dffe_12,
	dffe2,
	dffe3,
	dffe4,
	dffe5,
	dffe6,
	dffe7,
	dffe8,
	dffe9,
	dffe121,
	pipeline_dffe_11,
	dffe111,
	pipeline_dffe_10,
	dffe91,
	dffe101,
	pipeline_dffe_8,
	pipeline_dffe_9,
	dffe19,
	dffe21,
	dffe31,
	dffe41,
	dffe51,
	dffe61,
	dffe71,
	dffe81,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	sin_o_0;
output 	dffe18;
output 	dffe17;
input 	dffe16;
input 	pipeline_dffe_17;
output 	dffe161;
input 	dffe181;
output 	dffe15;
input 	dffe171;
output 	dffe14;
input 	pipeline_dffe_16;
input 	dffe162;
output 	dffe13;
input 	pipeline_dffe_15;
input 	dffe151;
output 	dffe12;
input 	pipeline_dffe_14;
output 	dffe10;
output 	dffe11;
input 	dffe141;
input 	pipeline_dffe_13;
input 	dffe131;
output 	dffe1;
input 	pipeline_dffe_12;
output 	dffe2;
output 	dffe3;
output 	dffe4;
output 	dffe5;
output 	dffe6;
output 	dffe7;
output 	dffe8;
output 	dffe9;
input 	dffe121;
input 	pipeline_dffe_11;
input 	dffe111;
input 	pipeline_dffe_10;
input 	dffe91;
input 	dffe101;
input 	pipeline_dffe_8;
input 	pipeline_dffe_9;
input 	dffe19;
input 	dffe21;
input 	dffe31;
input 	dffe41;
input 	dffe51;
input 	dffe61;
input 	dffe71;
input 	dffe81;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[17]~q ;
wire \xordvalue[10]~q ;
wire \Add0~1_sumout ;
wire \a[16]~q ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \a[15]~q ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \a[14]~q ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \a[13]~q ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \a[12]~q ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \a[11]~q ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \a[10]~q ;
wire \a[9]~q ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \a[8]~q ;
wire \xordvalue[8]~q ;
wire \a[0]~q ;
wire \xordvalue[0]~q ;
wire \a[1]~q ;
wire \xordvalue[1]~q ;
wire \a[2]~q ;
wire \xordvalue[2]~q ;
wire \a[3]~q ;
wire \xordvalue[3]~q ;
wire \a[4]~q ;
wire \xordvalue[4]~q ;
wire \a[5]~q ;
wire \xordvalue[5]~q ;
wire \a[6]~q ;
wire \xordvalue[6]~q ;
wire \a[7]~q ;
wire \xordvalue[7]~q ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~51 ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~55 ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~59 ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~63 ;
wire \Add0~65_sumout ;
wire \Add0~66 ;
wire \Add0~67 ;
wire \Add0~69_sumout ;
wire \Add0~70 ;
wire \Add0~71 ;
wire \xordvalue~0_combout ;
wire \xordvalue~1_combout ;
wire \xordvalue~2_combout ;
wire \xordvalue~3_combout ;
wire \xordvalue~4_combout ;
wire \xordvalue~5_combout ;
wire \xordvalue~6_combout ;
wire \xordvalue~7_combout ;
wire \xordvalue~8_combout ;
wire \xordvalue~9_combout ;


nco_test_lpm_add_sub_24 u0(
	.a_17(\a[17]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.a_16(\a[16]~q ),
	.a_15(\a[15]~q ),
	.a_14(\a[14]~q ),
	.a_13(\a[13]~q ),
	.a_12(\a[12]~q ),
	.a_11(\a[11]~q ),
	.a_10(\a[10]~q ),
	.a_9(\a[9]~q ),
	.a_8(\a[8]~q ),
	.xordvalue_8(\xordvalue[8]~q ),
	.a_0(\a[0]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_1(\a[1]~q ),
	.xordvalue_1(\xordvalue[1]~q ),
	.a_2(\a[2]~q ),
	.xordvalue_2(\xordvalue[2]~q ),
	.a_3(\a[3]~q ),
	.xordvalue_3(\xordvalue[3]~q ),
	.a_4(\a[4]~q ),
	.xordvalue_4(\xordvalue[4]~q ),
	.a_5(\a[5]~q ),
	.xordvalue_5(\xordvalue[5]~q ),
	.a_6(\a[6]~q ),
	.xordvalue_6(\xordvalue[6]~q ),
	.a_7(\a[7]~q ),
	.xordvalue_7(\xordvalue[7]~q ),
	.dffe18(dffe18),
	.dffe17(dffe17),
	.dffe16(dffe161),
	.dffe15(dffe15),
	.dffe14(dffe14),
	.dffe13(dffe13),
	.dffe12(dffe12),
	.dffe10(dffe10),
	.dffe11(dffe11),
	.dffe1(dffe1),
	.dffe2(dffe2),
	.dffe3(dffe3),
	.dffe4(dffe4),
	.dffe5(dffe5),
	.dffe6(dffe6),
	.dffe7(dffe7),
	.dffe8(dffe8),
	.dffe9(dffe9),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[17] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[17]~q ),
	.prn(vcc));
defparam \a[17] .is_wysiwyg = "true";
defparam \a[17] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe181),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "on";

dffeas \a[16] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[16]~q ),
	.prn(vcc));
defparam \a[16] .is_wysiwyg = "true";
defparam \a[16] .power_up = "low";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe171),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~5 .shared_arith = "on";

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe162),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~9 .shared_arith = "on";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~13 .shared_arith = "on";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~17 .shared_arith = "on";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "on";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~25 .shared_arith = "on";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~29 .shared_arith = "on";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~33 .shared_arith = "on";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \xordvalue[8] (
	.clk(clk),
	.d(\xordvalue~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[8]~q ),
	.prn(vcc));
defparam \xordvalue[8] .is_wysiwyg = "true";
defparam \xordvalue[8] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \xordvalue[1] (
	.clk(clk),
	.d(\xordvalue~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[1]~q ),
	.prn(vcc));
defparam \xordvalue[1] .is_wysiwyg = "true";
defparam \xordvalue[1] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \xordvalue[2] (
	.clk(clk),
	.d(\xordvalue~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[2]~q ),
	.prn(vcc));
defparam \xordvalue[2] .is_wysiwyg = "true";
defparam \xordvalue[2] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \xordvalue[3] (
	.clk(clk),
	.d(\xordvalue~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[3]~q ),
	.prn(vcc));
defparam \xordvalue[3] .is_wysiwyg = "true";
defparam \xordvalue[3] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \xordvalue[4] (
	.clk(clk),
	.d(\xordvalue~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[4]~q ),
	.prn(vcc));
defparam \xordvalue[4] .is_wysiwyg = "true";
defparam \xordvalue[4] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \xordvalue[5] (
	.clk(clk),
	.d(\xordvalue~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[5]~q ),
	.prn(vcc));
defparam \xordvalue[5] .is_wysiwyg = "true";
defparam \xordvalue[5] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \xordvalue[6] (
	.clk(clk),
	.d(\xordvalue~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[6]~q ),
	.prn(vcc));
defparam \xordvalue[6] .is_wysiwyg = "true";
defparam \xordvalue[6] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \xordvalue[7] (
	.clk(clk),
	.d(\xordvalue~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[7]~q ),
	.prn(vcc));
defparam \xordvalue[7] .is_wysiwyg = "true";
defparam \xordvalue[7] .power_up = "low";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~70 ),
	.sharein(\Add0~71 ),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~37 .shared_arith = "on";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!dffe19),
	.datad(!dffe16),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add0~41 .shared_arith = "on";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout(\Add0~47 ));
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~45 .shared_arith = "on";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(\Add0~47 ),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout(\Add0~51 ));
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~49 .shared_arith = "on";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(\Add0~51 ),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout(\Add0~55 ));
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~53 .shared_arith = "on";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(\Add0~55 ),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout(\Add0~59 ));
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~57 .shared_arith = "on";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(\Add0~59 ),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout(\Add0~63 ));
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~61 .shared_arith = "on";

arriav_lcell_comb \Add0~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(\Add0~63 ),
	.combout(),
	.sumout(\Add0~65_sumout ),
	.cout(\Add0~66 ),
	.shareout(\Add0~67 ));
defparam \Add0~65 .extended_lut = "off";
defparam \Add0~65 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~65 .shared_arith = "on";

arriav_lcell_comb \Add0~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~66 ),
	.sharein(\Add0~67 ),
	.combout(),
	.sumout(\Add0~69_sumout ),
	.cout(\Add0~70 ),
	.shareout(\Add0~71 ));
defparam \Add0~69 .extended_lut = "off";
defparam \Add0~69 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~69 .shared_arith = "on";

arriav_lcell_comb \xordvalue~0 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_17),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

arriav_lcell_comb \xordvalue~1 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~1 .extended_lut = "off";
defparam \xordvalue~1 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~1 .shared_arith = "off";

arriav_lcell_comb \xordvalue~2 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_8),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~2 .extended_lut = "off";
defparam \xordvalue~2 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~2 .shared_arith = "off";

arriav_lcell_comb \xordvalue~3 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_9),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~3 .extended_lut = "off";
defparam \xordvalue~3 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~3 .shared_arith = "off";

arriav_lcell_comb \xordvalue~4 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_10),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~4 .extended_lut = "off";
defparam \xordvalue~4 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~4 .shared_arith = "off";

arriav_lcell_comb \xordvalue~5 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_11),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~5 .extended_lut = "off";
defparam \xordvalue~5 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~5 .shared_arith = "off";

arriav_lcell_comb \xordvalue~6 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_12),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~6 .extended_lut = "off";
defparam \xordvalue~6 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~6 .shared_arith = "off";

arriav_lcell_comb \xordvalue~7 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_13),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~7 .extended_lut = "off";
defparam \xordvalue~7 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~7 .shared_arith = "off";

arriav_lcell_comb \xordvalue~8 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_14),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~8 .extended_lut = "off";
defparam \xordvalue~8 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~8 .shared_arith = "off";

arriav_lcell_comb \xordvalue~9 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_15),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~9 .extended_lut = "off";
defparam \xordvalue~9 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~9 .shared_arith = "off";

endmodule

module nco_test_lpm_add_sub_24 (
	a_17,
	xordvalue_10,
	a_16,
	a_15,
	a_14,
	a_13,
	a_12,
	a_11,
	a_10,
	a_9,
	a_8,
	xordvalue_8,
	a_0,
	xordvalue_0,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	a_4,
	xordvalue_4,
	a_5,
	xordvalue_5,
	a_6,
	xordvalue_6,
	a_7,
	xordvalue_7,
	dffe18,
	dffe17,
	dffe16,
	dffe15,
	dffe14,
	dffe13,
	dffe12,
	dffe10,
	dffe11,
	dffe1,
	dffe2,
	dffe3,
	dffe4,
	dffe5,
	dffe6,
	dffe7,
	dffe8,
	dffe9,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_10;
input 	a_16;
input 	a_15;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_10;
input 	a_9;
input 	a_8;
input 	xordvalue_8;
input 	a_0;
input 	xordvalue_0;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
input 	a_4;
input 	xordvalue_4;
input 	a_5;
input 	xordvalue_5;
input 	a_6;
input 	xordvalue_6;
input 	a_7;
input 	xordvalue_7;
output 	dffe18;
output 	dffe17;
output 	dffe16;
output 	dffe15;
output 	dffe14;
output 	dffe13;
output 	dffe12;
output 	dffe10;
output 	dffe11;
output 	dffe1;
output 	dffe2;
output 	dffe3;
output 	dffe4;
output 	dffe5;
output 	dffe6;
output 	dffe7;
output 	dffe8;
output 	dffe9;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_add_sub_jdg_5 auto_generated(
	.a_17(a_17),
	.xordvalue_10(xordvalue_10),
	.a_16(a_16),
	.a_15(a_15),
	.a_14(a_14),
	.a_13(a_13),
	.a_12(a_12),
	.a_11(a_11),
	.a_10(a_10),
	.a_9(a_9),
	.a_8(a_8),
	.xordvalue_8(xordvalue_8),
	.a_0(a_0),
	.xordvalue_0(xordvalue_0),
	.a_1(a_1),
	.xordvalue_1(xordvalue_1),
	.a_2(a_2),
	.xordvalue_2(xordvalue_2),
	.a_3(a_3),
	.xordvalue_3(xordvalue_3),
	.a_4(a_4),
	.xordvalue_4(xordvalue_4),
	.a_5(a_5),
	.xordvalue_5(xordvalue_5),
	.a_6(a_6),
	.xordvalue_6(xordvalue_6),
	.a_7(a_7),
	.xordvalue_7(xordvalue_7),
	.dffe181(dffe18),
	.dffe171(dffe17),
	.dffe161(dffe16),
	.dffe151(dffe15),
	.dffe141(dffe14),
	.dffe131(dffe13),
	.dffe121(dffe12),
	.dffe101(dffe10),
	.dffe111(dffe11),
	.dffe19(dffe1),
	.dffe21(dffe2),
	.dffe31(dffe3),
	.dffe41(dffe4),
	.dffe51(dffe5),
	.dffe61(dffe6),
	.dffe71(dffe7),
	.dffe81(dffe8),
	.dffe91(dffe9),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module nco_test_add_sub_jdg_5 (
	a_17,
	xordvalue_10,
	a_16,
	a_15,
	a_14,
	a_13,
	a_12,
	a_11,
	a_10,
	a_9,
	a_8,
	xordvalue_8,
	a_0,
	xordvalue_0,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	a_4,
	xordvalue_4,
	a_5,
	xordvalue_5,
	a_6,
	xordvalue_6,
	a_7,
	xordvalue_7,
	dffe181,
	dffe171,
	dffe161,
	dffe151,
	dffe141,
	dffe131,
	dffe121,
	dffe101,
	dffe111,
	dffe19,
	dffe21,
	dffe31,
	dffe41,
	dffe51,
	dffe61,
	dffe71,
	dffe81,
	dffe91,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_10;
input 	a_16;
input 	a_15;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_10;
input 	a_9;
input 	a_8;
input 	xordvalue_8;
input 	a_0;
input 	xordvalue_0;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
input 	a_4;
input 	xordvalue_4;
input 	a_5;
input 	xordvalue_5;
input 	a_6;
input 	xordvalue_6;
input 	a_7;
input 	xordvalue_7;
output 	dffe181;
output 	dffe171;
output 	dffe161;
output 	dffe151;
output 	dffe141;
output 	dffe131;
output 	dffe121;
output 	dffe101;
output 	dffe111;
output 	dffe19;
output 	dffe21;
output 	dffe31;
output 	dffe41;
output 	dffe51;
output 	dffe61;
output 	dffe71;
output 	dffe81;
output 	dffe91;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~COUT ;
wire \add_sub_cella[12]~COUT ;
wire \add_sub_cella[13]~COUT ;
wire \add_sub_cella[14]~COUT ;
wire \add_sub_cella[15]~COUT ;
wire \add_sub_cella[16]~COUT ;
wire \add_sub_cella[17]~sumout ;
wire \add_sub_cella[16]~sumout ;
wire \add_sub_cella[15]~sumout ;
wire \add_sub_cella[14]~sumout ;
wire \add_sub_cella[13]~sumout ;
wire \add_sub_cella[12]~sumout ;
wire \add_sub_cella[11]~sumout ;
wire \add_sub_cella[9]~sumout ;
wire \add_sub_cella[10]~sumout ;
wire \add_sub_cella[0]~sumout ;
wire \add_sub_cella[1]~sumout ;
wire \add_sub_cella[2]~sumout ;
wire \add_sub_cella[3]~sumout ;
wire \add_sub_cella[4]~sumout ;
wire \add_sub_cella[5]~sumout ;
wire \add_sub_cella[6]~sumout ;
wire \add_sub_cella[7]~sumout ;
wire \add_sub_cella[8]~sumout ;


dffeas dffe18(
	.clk(clock),
	.d(\add_sub_cella[17]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe181),
	.prn(vcc));
defparam dffe18.is_wysiwyg = "true";
defparam dffe18.power_up = "low";

dffeas dffe17(
	.clk(clock),
	.d(\add_sub_cella[16]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe171),
	.prn(vcc));
defparam dffe17.is_wysiwyg = "true";
defparam dffe17.power_up = "low";

dffeas dffe16(
	.clk(clock),
	.d(\add_sub_cella[15]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe161),
	.prn(vcc));
defparam dffe16.is_wysiwyg = "true";
defparam dffe16.power_up = "low";

dffeas dffe15(
	.clk(clock),
	.d(\add_sub_cella[14]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe151),
	.prn(vcc));
defparam dffe15.is_wysiwyg = "true";
defparam dffe15.power_up = "low";

dffeas dffe14(
	.clk(clock),
	.d(\add_sub_cella[13]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe141),
	.prn(vcc));
defparam dffe14.is_wysiwyg = "true";
defparam dffe14.power_up = "low";

dffeas dffe13(
	.clk(clock),
	.d(\add_sub_cella[12]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe131),
	.prn(vcc));
defparam dffe13.is_wysiwyg = "true";
defparam dffe13.power_up = "low";

dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe19),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

arriav_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_1),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_2),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_3),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_4),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_5),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_6),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_7),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_8),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(\add_sub_cella[11]~COUT ),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[12] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[11]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[12]~sumout ),
	.cout(\add_sub_cella[12]~COUT ),
	.shareout());
defparam \add_sub_cella[12] .extended_lut = "off";
defparam \add_sub_cella[12] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[12] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[13] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[12]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[13]~sumout ),
	.cout(\add_sub_cella[13]~COUT ),
	.shareout());
defparam \add_sub_cella[13] .extended_lut = "off";
defparam \add_sub_cella[13] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[13] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[14] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[13]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[14]~sumout ),
	.cout(\add_sub_cella[14]~COUT ),
	.shareout());
defparam \add_sub_cella[14] .extended_lut = "off";
defparam \add_sub_cella[14] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[14] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[15] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[14]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[15]~sumout ),
	.cout(\add_sub_cella[15]~COUT ),
	.shareout());
defparam \add_sub_cella[15] .extended_lut = "off";
defparam \add_sub_cella[15] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[15] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[16] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_16),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[15]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[16]~sumout ),
	.cout(\add_sub_cella[16]~COUT ),
	.shareout());
defparam \add_sub_cella[16] .extended_lut = "off";
defparam \add_sub_cella[16] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[16] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[17] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_17),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[16]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[17]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[17] .extended_lut = "off";
defparam \add_sub_cella[17] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[17] .shared_arith = "off";

endmodule

module nco_test_cordic_sxor_1p_lpm_6 (
	sin_o_0,
	dffe18,
	dffe17,
	dffe16,
	dffe161,
	dffe181,
	pipeline_dffe_17,
	dffe15,
	dffe14,
	pipeline_dffe_16,
	dffe171,
	dffe13,
	pipeline_dffe_15,
	dffe162,
	dffe11,
	dffe12,
	pipeline_dffe_14,
	dffe151,
	pipeline_dffe_13,
	dffe1,
	dffe141,
	dffe2,
	dffe3,
	dffe4,
	dffe5,
	dffe6,
	dffe7,
	dffe8,
	dffe9,
	dffe10,
	pipeline_dffe_12,
	dffe131,
	pipeline_dffe_11,
	dffe121,
	dffe101,
	dffe111,
	pipeline_dffe_10,
	pipeline_dffe_9,
	dffe19,
	dffe21,
	dffe31,
	dffe41,
	dffe51,
	dffe61,
	dffe71,
	dffe81,
	dffe91,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	sin_o_0;
output 	dffe18;
output 	dffe17;
input 	dffe16;
output 	dffe161;
input 	dffe181;
input 	pipeline_dffe_17;
output 	dffe15;
output 	dffe14;
input 	pipeline_dffe_16;
input 	dffe171;
output 	dffe13;
input 	pipeline_dffe_15;
input 	dffe162;
output 	dffe11;
output 	dffe12;
input 	pipeline_dffe_14;
input 	dffe151;
input 	pipeline_dffe_13;
output 	dffe1;
input 	dffe141;
output 	dffe2;
output 	dffe3;
output 	dffe4;
output 	dffe5;
output 	dffe6;
output 	dffe7;
output 	dffe8;
output 	dffe9;
output 	dffe10;
input 	pipeline_dffe_12;
input 	dffe131;
input 	pipeline_dffe_11;
input 	dffe121;
input 	dffe101;
input 	dffe111;
input 	pipeline_dffe_10;
input 	pipeline_dffe_9;
input 	dffe19;
input 	dffe21;
input 	dffe31;
input 	dffe41;
input 	dffe51;
input 	dffe61;
input 	dffe71;
input 	dffe81;
input 	dffe91;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[17]~q ;
wire \xordvalue[10]~q ;
wire \Add0~1_sumout ;
wire \a[16]~q ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \a[15]~q ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \a[14]~q ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \a[13]~q ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \a[12]~q ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \a[11]~q ;
wire \a[10]~q ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \a[9]~q ;
wire \a[0]~q ;
wire \xordvalue[0]~q ;
wire \a[1]~q ;
wire \xordvalue[1]~q ;
wire \a[2]~q ;
wire \xordvalue[2]~q ;
wire \a[3]~q ;
wire \xordvalue[3]~q ;
wire \a[4]~q ;
wire \xordvalue[4]~q ;
wire \a[5]~q ;
wire \xordvalue[5]~q ;
wire \a[6]~q ;
wire \xordvalue[6]~q ;
wire \a[7]~q ;
wire \xordvalue[7]~q ;
wire \a[8]~q ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~51 ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~55 ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~59 ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~63 ;
wire \Add0~65_sumout ;
wire \Add0~66 ;
wire \Add0~67 ;
wire \Add0~69_sumout ;
wire \Add0~70 ;
wire \Add0~71 ;
wire \xordvalue~0_combout ;
wire \xordvalue~1_combout ;
wire \xordvalue~2_combout ;
wire \xordvalue~3_combout ;
wire \xordvalue~4_combout ;
wire \xordvalue~5_combout ;
wire \xordvalue~6_combout ;
wire \xordvalue~7_combout ;
wire \xordvalue~8_combout ;


nco_test_lpm_add_sub_25 u0(
	.a_17(\a[17]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.a_16(\a[16]~q ),
	.a_15(\a[15]~q ),
	.a_14(\a[14]~q ),
	.a_13(\a[13]~q ),
	.a_12(\a[12]~q ),
	.a_11(\a[11]~q ),
	.a_10(\a[10]~q ),
	.a_9(\a[9]~q ),
	.a_0(\a[0]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_1(\a[1]~q ),
	.xordvalue_1(\xordvalue[1]~q ),
	.a_2(\a[2]~q ),
	.xordvalue_2(\xordvalue[2]~q ),
	.a_3(\a[3]~q ),
	.xordvalue_3(\xordvalue[3]~q ),
	.a_4(\a[4]~q ),
	.xordvalue_4(\xordvalue[4]~q ),
	.a_5(\a[5]~q ),
	.xordvalue_5(\xordvalue[5]~q ),
	.a_6(\a[6]~q ),
	.xordvalue_6(\xordvalue[6]~q ),
	.a_7(\a[7]~q ),
	.xordvalue_7(\xordvalue[7]~q ),
	.a_8(\a[8]~q ),
	.dffe18(dffe18),
	.dffe17(dffe17),
	.dffe16(dffe161),
	.dffe15(dffe15),
	.dffe14(dffe14),
	.dffe13(dffe13),
	.dffe11(dffe11),
	.dffe12(dffe12),
	.dffe1(dffe1),
	.dffe2(dffe2),
	.dffe3(dffe3),
	.dffe4(dffe4),
	.dffe5(dffe5),
	.dffe6(dffe6),
	.dffe7(dffe7),
	.dffe8(dffe8),
	.dffe9(dffe9),
	.dffe10(dffe10),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[17] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[17]~q ),
	.prn(vcc));
defparam \a[17] .is_wysiwyg = "true";
defparam \a[17] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe181),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "on";

dffeas \a[16] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[16]~q ),
	.prn(vcc));
defparam \a[16] .is_wysiwyg = "true";
defparam \a[16] .power_up = "low";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe171),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~5 .shared_arith = "on";

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe162),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~9 .shared_arith = "on";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~13 .shared_arith = "on";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~17 .shared_arith = "on";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "on";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~25 .shared_arith = "on";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~29 .shared_arith = "on";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \xordvalue[1] (
	.clk(clk),
	.d(\xordvalue~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[1]~q ),
	.prn(vcc));
defparam \xordvalue[1] .is_wysiwyg = "true";
defparam \xordvalue[1] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \xordvalue[2] (
	.clk(clk),
	.d(\xordvalue~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[2]~q ),
	.prn(vcc));
defparam \xordvalue[2] .is_wysiwyg = "true";
defparam \xordvalue[2] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \xordvalue[3] (
	.clk(clk),
	.d(\xordvalue~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[3]~q ),
	.prn(vcc));
defparam \xordvalue[3] .is_wysiwyg = "true";
defparam \xordvalue[3] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \xordvalue[4] (
	.clk(clk),
	.d(\xordvalue~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[4]~q ),
	.prn(vcc));
defparam \xordvalue[4] .is_wysiwyg = "true";
defparam \xordvalue[4] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \xordvalue[5] (
	.clk(clk),
	.d(\xordvalue~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[5]~q ),
	.prn(vcc));
defparam \xordvalue[5] .is_wysiwyg = "true";
defparam \xordvalue[5] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \xordvalue[6] (
	.clk(clk),
	.d(\xordvalue~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[6]~q ),
	.prn(vcc));
defparam \xordvalue[6] .is_wysiwyg = "true";
defparam \xordvalue[6] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \xordvalue[7] (
	.clk(clk),
	.d(\xordvalue~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[7]~q ),
	.prn(vcc));
defparam \xordvalue[7] .is_wysiwyg = "true";
defparam \xordvalue[7] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~70 ),
	.sharein(\Add0~71 ),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~33 .shared_arith = "on";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!dffe19),
	.datad(!dffe16),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add0~37 .shared_arith = "on";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~41 .shared_arith = "on";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout(\Add0~47 ));
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~45 .shared_arith = "on";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(\Add0~47 ),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout(\Add0~51 ));
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~49 .shared_arith = "on";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(\Add0~51 ),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout(\Add0~55 ));
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~53 .shared_arith = "on";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(\Add0~55 ),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout(\Add0~59 ));
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~57 .shared_arith = "on";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(\Add0~59 ),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout(\Add0~63 ));
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~61 .shared_arith = "on";

arriav_lcell_comb \Add0~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(\Add0~63 ),
	.combout(),
	.sumout(\Add0~65_sumout ),
	.cout(\Add0~66 ),
	.shareout(\Add0~67 ));
defparam \Add0~65 .extended_lut = "off";
defparam \Add0~65 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~65 .shared_arith = "on";

arriav_lcell_comb \Add0~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~66 ),
	.sharein(\Add0~67 ),
	.combout(),
	.sumout(\Add0~69_sumout ),
	.cout(\Add0~70 ),
	.shareout(\Add0~71 ));
defparam \Add0~69 .extended_lut = "off";
defparam \Add0~69 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~69 .shared_arith = "on";

arriav_lcell_comb \xordvalue~0 (
	.dataa(!pipeline_dffe_17),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

arriav_lcell_comb \xordvalue~1 (
	.dataa(!pipeline_dffe_9),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~1 .extended_lut = "off";
defparam \xordvalue~1 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~1 .shared_arith = "off";

arriav_lcell_comb \xordvalue~2 (
	.dataa(!pipeline_dffe_10),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~2 .extended_lut = "off";
defparam \xordvalue~2 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~2 .shared_arith = "off";

arriav_lcell_comb \xordvalue~3 (
	.dataa(!pipeline_dffe_11),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~3 .extended_lut = "off";
defparam \xordvalue~3 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~3 .shared_arith = "off";

arriav_lcell_comb \xordvalue~4 (
	.dataa(!pipeline_dffe_12),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~4 .extended_lut = "off";
defparam \xordvalue~4 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~4 .shared_arith = "off";

arriav_lcell_comb \xordvalue~5 (
	.dataa(!pipeline_dffe_13),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~5 .extended_lut = "off";
defparam \xordvalue~5 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~5 .shared_arith = "off";

arriav_lcell_comb \xordvalue~6 (
	.dataa(!pipeline_dffe_14),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~6 .extended_lut = "off";
defparam \xordvalue~6 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~6 .shared_arith = "off";

arriav_lcell_comb \xordvalue~7 (
	.dataa(!pipeline_dffe_15),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~7 .extended_lut = "off";
defparam \xordvalue~7 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~7 .shared_arith = "off";

arriav_lcell_comb \xordvalue~8 (
	.dataa(!pipeline_dffe_16),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~8 .extended_lut = "off";
defparam \xordvalue~8 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~8 .shared_arith = "off";

endmodule

module nco_test_lpm_add_sub_25 (
	a_17,
	xordvalue_10,
	a_16,
	a_15,
	a_14,
	a_13,
	a_12,
	a_11,
	a_10,
	a_9,
	a_0,
	xordvalue_0,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	a_4,
	xordvalue_4,
	a_5,
	xordvalue_5,
	a_6,
	xordvalue_6,
	a_7,
	xordvalue_7,
	a_8,
	dffe18,
	dffe17,
	dffe16,
	dffe15,
	dffe14,
	dffe13,
	dffe11,
	dffe12,
	dffe1,
	dffe2,
	dffe3,
	dffe4,
	dffe5,
	dffe6,
	dffe7,
	dffe8,
	dffe9,
	dffe10,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_10;
input 	a_16;
input 	a_15;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_10;
input 	a_9;
input 	a_0;
input 	xordvalue_0;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
input 	a_4;
input 	xordvalue_4;
input 	a_5;
input 	xordvalue_5;
input 	a_6;
input 	xordvalue_6;
input 	a_7;
input 	xordvalue_7;
input 	a_8;
output 	dffe18;
output 	dffe17;
output 	dffe16;
output 	dffe15;
output 	dffe14;
output 	dffe13;
output 	dffe11;
output 	dffe12;
output 	dffe1;
output 	dffe2;
output 	dffe3;
output 	dffe4;
output 	dffe5;
output 	dffe6;
output 	dffe7;
output 	dffe8;
output 	dffe9;
output 	dffe10;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_add_sub_jdg_6 auto_generated(
	.a_17(a_17),
	.xordvalue_10(xordvalue_10),
	.a_16(a_16),
	.a_15(a_15),
	.a_14(a_14),
	.a_13(a_13),
	.a_12(a_12),
	.a_11(a_11),
	.a_10(a_10),
	.a_9(a_9),
	.a_0(a_0),
	.xordvalue_0(xordvalue_0),
	.a_1(a_1),
	.xordvalue_1(xordvalue_1),
	.a_2(a_2),
	.xordvalue_2(xordvalue_2),
	.a_3(a_3),
	.xordvalue_3(xordvalue_3),
	.a_4(a_4),
	.xordvalue_4(xordvalue_4),
	.a_5(a_5),
	.xordvalue_5(xordvalue_5),
	.a_6(a_6),
	.xordvalue_6(xordvalue_6),
	.a_7(a_7),
	.xordvalue_7(xordvalue_7),
	.a_8(a_8),
	.dffe181(dffe18),
	.dffe171(dffe17),
	.dffe161(dffe16),
	.dffe151(dffe15),
	.dffe141(dffe14),
	.dffe131(dffe13),
	.dffe111(dffe11),
	.dffe121(dffe12),
	.dffe19(dffe1),
	.dffe21(dffe2),
	.dffe31(dffe3),
	.dffe41(dffe4),
	.dffe51(dffe5),
	.dffe61(dffe6),
	.dffe71(dffe7),
	.dffe81(dffe8),
	.dffe91(dffe9),
	.dffe101(dffe10),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module nco_test_add_sub_jdg_6 (
	a_17,
	xordvalue_10,
	a_16,
	a_15,
	a_14,
	a_13,
	a_12,
	a_11,
	a_10,
	a_9,
	a_0,
	xordvalue_0,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	a_4,
	xordvalue_4,
	a_5,
	xordvalue_5,
	a_6,
	xordvalue_6,
	a_7,
	xordvalue_7,
	a_8,
	dffe181,
	dffe171,
	dffe161,
	dffe151,
	dffe141,
	dffe131,
	dffe111,
	dffe121,
	dffe19,
	dffe21,
	dffe31,
	dffe41,
	dffe51,
	dffe61,
	dffe71,
	dffe81,
	dffe91,
	dffe101,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_10;
input 	a_16;
input 	a_15;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_10;
input 	a_9;
input 	a_0;
input 	xordvalue_0;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
input 	a_4;
input 	xordvalue_4;
input 	a_5;
input 	xordvalue_5;
input 	a_6;
input 	xordvalue_6;
input 	a_7;
input 	xordvalue_7;
input 	a_8;
output 	dffe181;
output 	dffe171;
output 	dffe161;
output 	dffe151;
output 	dffe141;
output 	dffe131;
output 	dffe111;
output 	dffe121;
output 	dffe19;
output 	dffe21;
output 	dffe31;
output 	dffe41;
output 	dffe51;
output 	dffe61;
output 	dffe71;
output 	dffe81;
output 	dffe91;
output 	dffe101;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~COUT ;
wire \add_sub_cella[12]~COUT ;
wire \add_sub_cella[13]~COUT ;
wire \add_sub_cella[14]~COUT ;
wire \add_sub_cella[15]~COUT ;
wire \add_sub_cella[16]~COUT ;
wire \add_sub_cella[17]~sumout ;
wire \add_sub_cella[16]~sumout ;
wire \add_sub_cella[15]~sumout ;
wire \add_sub_cella[14]~sumout ;
wire \add_sub_cella[13]~sumout ;
wire \add_sub_cella[12]~sumout ;
wire \add_sub_cella[10]~sumout ;
wire \add_sub_cella[11]~sumout ;
wire \add_sub_cella[0]~sumout ;
wire \add_sub_cella[1]~sumout ;
wire \add_sub_cella[2]~sumout ;
wire \add_sub_cella[3]~sumout ;
wire \add_sub_cella[4]~sumout ;
wire \add_sub_cella[5]~sumout ;
wire \add_sub_cella[6]~sumout ;
wire \add_sub_cella[7]~sumout ;
wire \add_sub_cella[8]~sumout ;
wire \add_sub_cella[9]~sumout ;


dffeas dffe18(
	.clk(clock),
	.d(\add_sub_cella[17]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe181),
	.prn(vcc));
defparam dffe18.is_wysiwyg = "true";
defparam dffe18.power_up = "low";

dffeas dffe17(
	.clk(clock),
	.d(\add_sub_cella[16]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe171),
	.prn(vcc));
defparam dffe17.is_wysiwyg = "true";
defparam dffe17.power_up = "low";

dffeas dffe16(
	.clk(clock),
	.d(\add_sub_cella[15]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe161),
	.prn(vcc));
defparam dffe16.is_wysiwyg = "true";
defparam dffe16.power_up = "low";

dffeas dffe15(
	.clk(clock),
	.d(\add_sub_cella[14]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe151),
	.prn(vcc));
defparam dffe15.is_wysiwyg = "true";
defparam dffe15.power_up = "low";

dffeas dffe14(
	.clk(clock),
	.d(\add_sub_cella[13]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe141),
	.prn(vcc));
defparam dffe14.is_wysiwyg = "true";
defparam dffe14.power_up = "low";

dffeas dffe13(
	.clk(clock),
	.d(\add_sub_cella[12]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe131),
	.prn(vcc));
defparam dffe13.is_wysiwyg = "true";
defparam dffe13.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe19),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

arriav_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_1),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_2),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_3),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_4),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_5),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_6),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_7),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(\add_sub_cella[11]~COUT ),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[12] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[11]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[12]~sumout ),
	.cout(\add_sub_cella[12]~COUT ),
	.shareout());
defparam \add_sub_cella[12] .extended_lut = "off";
defparam \add_sub_cella[12] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[12] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[13] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[12]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[13]~sumout ),
	.cout(\add_sub_cella[13]~COUT ),
	.shareout());
defparam \add_sub_cella[13] .extended_lut = "off";
defparam \add_sub_cella[13] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[13] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[14] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[13]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[14]~sumout ),
	.cout(\add_sub_cella[14]~COUT ),
	.shareout());
defparam \add_sub_cella[14] .extended_lut = "off";
defparam \add_sub_cella[14] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[14] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[15] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[14]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[15]~sumout ),
	.cout(\add_sub_cella[15]~COUT ),
	.shareout());
defparam \add_sub_cella[15] .extended_lut = "off";
defparam \add_sub_cella[15] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[15] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[16] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_16),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[15]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[16]~sumout ),
	.cout(\add_sub_cella[16]~COUT ),
	.shareout());
defparam \add_sub_cella[16] .extended_lut = "off";
defparam \add_sub_cella[16] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[16] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[17] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_17),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[16]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[17]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[17] .extended_lut = "off";
defparam \add_sub_cella[17] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[17] .shared_arith = "off";

endmodule

module nco_test_cordic_sxor_1p_lpm_7 (
	sin_o_0,
	dffe18,
	dffe17,
	dffe16,
	pipeline_dffe_17,
	dffe161,
	dffe181,
	dffe15,
	dffe171,
	dffe14,
	pipeline_dffe_16,
	dffe12,
	dffe13,
	dffe162,
	pipeline_dffe_15,
	dffe151,
	dffe1,
	pipeline_dffe_14,
	dffe2,
	dffe3,
	dffe4,
	dffe5,
	dffe6,
	dffe7,
	dffe8,
	dffe9,
	dffe10,
	dffe11,
	dffe141,
	pipeline_dffe_13,
	dffe131,
	pipeline_dffe_12,
	dffe111,
	dffe121,
	pipeline_dffe_10,
	pipeline_dffe_11,
	dffe19,
	dffe21,
	dffe31,
	dffe41,
	dffe51,
	dffe61,
	dffe71,
	dffe81,
	dffe91,
	dffe101,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	sin_o_0;
output 	dffe18;
output 	dffe17;
input 	dffe16;
input 	pipeline_dffe_17;
output 	dffe161;
input 	dffe181;
output 	dffe15;
input 	dffe171;
output 	dffe14;
input 	pipeline_dffe_16;
output 	dffe12;
output 	dffe13;
input 	dffe162;
input 	pipeline_dffe_15;
input 	dffe151;
output 	dffe1;
input 	pipeline_dffe_14;
output 	dffe2;
output 	dffe3;
output 	dffe4;
output 	dffe5;
output 	dffe6;
output 	dffe7;
output 	dffe8;
output 	dffe9;
output 	dffe10;
output 	dffe11;
input 	dffe141;
input 	pipeline_dffe_13;
input 	dffe131;
input 	pipeline_dffe_12;
input 	dffe111;
input 	dffe121;
input 	pipeline_dffe_10;
input 	pipeline_dffe_11;
input 	dffe19;
input 	dffe21;
input 	dffe31;
input 	dffe41;
input 	dffe51;
input 	dffe61;
input 	dffe71;
input 	dffe81;
input 	dffe91;
input 	dffe101;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[17]~q ;
wire \xordvalue[10]~q ;
wire \Add0~1_sumout ;
wire \a[16]~q ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \a[15]~q ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \a[14]~q ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \a[13]~q ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \a[12]~q ;
wire \a[11]~q ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \a[10]~q ;
wire \a[0]~q ;
wire \xordvalue[0]~q ;
wire \a[1]~q ;
wire \xordvalue[1]~q ;
wire \a[2]~q ;
wire \xordvalue[2]~q ;
wire \a[3]~q ;
wire \xordvalue[3]~q ;
wire \a[4]~q ;
wire \xordvalue[4]~q ;
wire \a[5]~q ;
wire \xordvalue[5]~q ;
wire \a[6]~q ;
wire \xordvalue[6]~q ;
wire \a[7]~q ;
wire \a[8]~q ;
wire \a[9]~q ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~51 ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~55 ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~59 ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~63 ;
wire \Add0~65_sumout ;
wire \Add0~66 ;
wire \Add0~67 ;
wire \Add0~69_sumout ;
wire \Add0~70 ;
wire \Add0~71 ;
wire \xordvalue~0_combout ;
wire \xordvalue~1_combout ;
wire \xordvalue~2_combout ;
wire \xordvalue~3_combout ;
wire \xordvalue~4_combout ;
wire \xordvalue~5_combout ;
wire \xordvalue~6_combout ;
wire \xordvalue~7_combout ;


nco_test_lpm_add_sub_26 u0(
	.a_17(\a[17]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.a_16(\a[16]~q ),
	.a_15(\a[15]~q ),
	.a_14(\a[14]~q ),
	.a_13(\a[13]~q ),
	.a_12(\a[12]~q ),
	.a_11(\a[11]~q ),
	.a_10(\a[10]~q ),
	.a_0(\a[0]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_1(\a[1]~q ),
	.xordvalue_1(\xordvalue[1]~q ),
	.a_2(\a[2]~q ),
	.xordvalue_2(\xordvalue[2]~q ),
	.a_3(\a[3]~q ),
	.xordvalue_3(\xordvalue[3]~q ),
	.a_4(\a[4]~q ),
	.xordvalue_4(\xordvalue[4]~q ),
	.a_5(\a[5]~q ),
	.xordvalue_5(\xordvalue[5]~q ),
	.a_6(\a[6]~q ),
	.xordvalue_6(\xordvalue[6]~q ),
	.a_7(\a[7]~q ),
	.a_8(\a[8]~q ),
	.a_9(\a[9]~q ),
	.dffe18(dffe18),
	.dffe17(dffe17),
	.dffe16(dffe161),
	.dffe15(dffe15),
	.dffe14(dffe14),
	.dffe12(dffe12),
	.dffe13(dffe13),
	.dffe1(dffe1),
	.dffe2(dffe2),
	.dffe3(dffe3),
	.dffe4(dffe4),
	.dffe5(dffe5),
	.dffe6(dffe6),
	.dffe7(dffe7),
	.dffe8(dffe8),
	.dffe9(dffe9),
	.dffe10(dffe10),
	.dffe11(dffe11),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[17] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[17]~q ),
	.prn(vcc));
defparam \a[17] .is_wysiwyg = "true";
defparam \a[17] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe181),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "on";

dffeas \a[16] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[16]~q ),
	.prn(vcc));
defparam \a[16] .is_wysiwyg = "true";
defparam \a[16] .power_up = "low";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe171),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~5 .shared_arith = "on";

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe162),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~9 .shared_arith = "on";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~13 .shared_arith = "on";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~17 .shared_arith = "on";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "on";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~25 .shared_arith = "on";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \xordvalue[1] (
	.clk(clk),
	.d(\xordvalue~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[1]~q ),
	.prn(vcc));
defparam \xordvalue[1] .is_wysiwyg = "true";
defparam \xordvalue[1] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \xordvalue[2] (
	.clk(clk),
	.d(\xordvalue~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[2]~q ),
	.prn(vcc));
defparam \xordvalue[2] .is_wysiwyg = "true";
defparam \xordvalue[2] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \xordvalue[3] (
	.clk(clk),
	.d(\xordvalue~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[3]~q ),
	.prn(vcc));
defparam \xordvalue[3] .is_wysiwyg = "true";
defparam \xordvalue[3] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \xordvalue[4] (
	.clk(clk),
	.d(\xordvalue~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[4]~q ),
	.prn(vcc));
defparam \xordvalue[4] .is_wysiwyg = "true";
defparam \xordvalue[4] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \xordvalue[5] (
	.clk(clk),
	.d(\xordvalue~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[5]~q ),
	.prn(vcc));
defparam \xordvalue[5] .is_wysiwyg = "true";
defparam \xordvalue[5] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \xordvalue[6] (
	.clk(clk),
	.d(\xordvalue~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[6]~q ),
	.prn(vcc));
defparam \xordvalue[6] .is_wysiwyg = "true";
defparam \xordvalue[6] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~70 ),
	.sharein(\Add0~71 ),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~29 .shared_arith = "on";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!dffe19),
	.datad(!dffe16),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add0~33 .shared_arith = "on";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~37 .shared_arith = "on";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~41 .shared_arith = "on";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout(\Add0~47 ));
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~45 .shared_arith = "on";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(\Add0~47 ),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout(\Add0~51 ));
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~49 .shared_arith = "on";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(\Add0~51 ),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout(\Add0~55 ));
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~53 .shared_arith = "on";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(\Add0~55 ),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout(\Add0~59 ));
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~57 .shared_arith = "on";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(\Add0~59 ),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout(\Add0~63 ));
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~61 .shared_arith = "on";

arriav_lcell_comb \Add0~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(\Add0~63 ),
	.combout(),
	.sumout(\Add0~65_sumout ),
	.cout(\Add0~66 ),
	.shareout(\Add0~67 ));
defparam \Add0~65 .extended_lut = "off";
defparam \Add0~65 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~65 .shared_arith = "on";

arriav_lcell_comb \Add0~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~66 ),
	.sharein(\Add0~67 ),
	.combout(),
	.sumout(\Add0~69_sumout ),
	.cout(\Add0~70 ),
	.shareout(\Add0~71 ));
defparam \Add0~69 .extended_lut = "off";
defparam \Add0~69 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~69 .shared_arith = "on";

arriav_lcell_comb \xordvalue~0 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_17),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

arriav_lcell_comb \xordvalue~1 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_10),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~1 .extended_lut = "off";
defparam \xordvalue~1 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~1 .shared_arith = "off";

arriav_lcell_comb \xordvalue~2 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_11),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~2 .extended_lut = "off";
defparam \xordvalue~2 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~2 .shared_arith = "off";

arriav_lcell_comb \xordvalue~3 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_12),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~3 .extended_lut = "off";
defparam \xordvalue~3 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~3 .shared_arith = "off";

arriav_lcell_comb \xordvalue~4 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_13),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~4 .extended_lut = "off";
defparam \xordvalue~4 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~4 .shared_arith = "off";

arriav_lcell_comb \xordvalue~5 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_14),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~5 .extended_lut = "off";
defparam \xordvalue~5 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~5 .shared_arith = "off";

arriav_lcell_comb \xordvalue~6 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_15),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~6 .extended_lut = "off";
defparam \xordvalue~6 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~6 .shared_arith = "off";

arriav_lcell_comb \xordvalue~7 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~7 .extended_lut = "off";
defparam \xordvalue~7 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~7 .shared_arith = "off";

endmodule

module nco_test_lpm_add_sub_26 (
	a_17,
	xordvalue_10,
	a_16,
	a_15,
	a_14,
	a_13,
	a_12,
	a_11,
	a_10,
	a_0,
	xordvalue_0,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	a_4,
	xordvalue_4,
	a_5,
	xordvalue_5,
	a_6,
	xordvalue_6,
	a_7,
	a_8,
	a_9,
	dffe18,
	dffe17,
	dffe16,
	dffe15,
	dffe14,
	dffe12,
	dffe13,
	dffe1,
	dffe2,
	dffe3,
	dffe4,
	dffe5,
	dffe6,
	dffe7,
	dffe8,
	dffe9,
	dffe10,
	dffe11,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_10;
input 	a_16;
input 	a_15;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_10;
input 	a_0;
input 	xordvalue_0;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
input 	a_4;
input 	xordvalue_4;
input 	a_5;
input 	xordvalue_5;
input 	a_6;
input 	xordvalue_6;
input 	a_7;
input 	a_8;
input 	a_9;
output 	dffe18;
output 	dffe17;
output 	dffe16;
output 	dffe15;
output 	dffe14;
output 	dffe12;
output 	dffe13;
output 	dffe1;
output 	dffe2;
output 	dffe3;
output 	dffe4;
output 	dffe5;
output 	dffe6;
output 	dffe7;
output 	dffe8;
output 	dffe9;
output 	dffe10;
output 	dffe11;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_add_sub_jdg_7 auto_generated(
	.a_17(a_17),
	.xordvalue_10(xordvalue_10),
	.a_16(a_16),
	.a_15(a_15),
	.a_14(a_14),
	.a_13(a_13),
	.a_12(a_12),
	.a_11(a_11),
	.a_10(a_10),
	.a_0(a_0),
	.xordvalue_0(xordvalue_0),
	.a_1(a_1),
	.xordvalue_1(xordvalue_1),
	.a_2(a_2),
	.xordvalue_2(xordvalue_2),
	.a_3(a_3),
	.xordvalue_3(xordvalue_3),
	.a_4(a_4),
	.xordvalue_4(xordvalue_4),
	.a_5(a_5),
	.xordvalue_5(xordvalue_5),
	.a_6(a_6),
	.xordvalue_6(xordvalue_6),
	.a_7(a_7),
	.a_8(a_8),
	.a_9(a_9),
	.dffe181(dffe18),
	.dffe171(dffe17),
	.dffe161(dffe16),
	.dffe151(dffe15),
	.dffe141(dffe14),
	.dffe121(dffe12),
	.dffe131(dffe13),
	.dffe19(dffe1),
	.dffe21(dffe2),
	.dffe31(dffe3),
	.dffe41(dffe4),
	.dffe51(dffe5),
	.dffe61(dffe6),
	.dffe71(dffe7),
	.dffe81(dffe8),
	.dffe91(dffe9),
	.dffe101(dffe10),
	.dffe111(dffe11),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module nco_test_add_sub_jdg_7 (
	a_17,
	xordvalue_10,
	a_16,
	a_15,
	a_14,
	a_13,
	a_12,
	a_11,
	a_10,
	a_0,
	xordvalue_0,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	a_4,
	xordvalue_4,
	a_5,
	xordvalue_5,
	a_6,
	xordvalue_6,
	a_7,
	a_8,
	a_9,
	dffe181,
	dffe171,
	dffe161,
	dffe151,
	dffe141,
	dffe121,
	dffe131,
	dffe19,
	dffe21,
	dffe31,
	dffe41,
	dffe51,
	dffe61,
	dffe71,
	dffe81,
	dffe91,
	dffe101,
	dffe111,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_10;
input 	a_16;
input 	a_15;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_10;
input 	a_0;
input 	xordvalue_0;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
input 	a_4;
input 	xordvalue_4;
input 	a_5;
input 	xordvalue_5;
input 	a_6;
input 	xordvalue_6;
input 	a_7;
input 	a_8;
input 	a_9;
output 	dffe181;
output 	dffe171;
output 	dffe161;
output 	dffe151;
output 	dffe141;
output 	dffe121;
output 	dffe131;
output 	dffe19;
output 	dffe21;
output 	dffe31;
output 	dffe41;
output 	dffe51;
output 	dffe61;
output 	dffe71;
output 	dffe81;
output 	dffe91;
output 	dffe101;
output 	dffe111;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~COUT ;
wire \add_sub_cella[12]~COUT ;
wire \add_sub_cella[13]~COUT ;
wire \add_sub_cella[14]~COUT ;
wire \add_sub_cella[15]~COUT ;
wire \add_sub_cella[16]~COUT ;
wire \add_sub_cella[17]~sumout ;
wire \add_sub_cella[16]~sumout ;
wire \add_sub_cella[15]~sumout ;
wire \add_sub_cella[14]~sumout ;
wire \add_sub_cella[13]~sumout ;
wire \add_sub_cella[11]~sumout ;
wire \add_sub_cella[12]~sumout ;
wire \add_sub_cella[0]~sumout ;
wire \add_sub_cella[1]~sumout ;
wire \add_sub_cella[2]~sumout ;
wire \add_sub_cella[3]~sumout ;
wire \add_sub_cella[4]~sumout ;
wire \add_sub_cella[5]~sumout ;
wire \add_sub_cella[6]~sumout ;
wire \add_sub_cella[7]~sumout ;
wire \add_sub_cella[8]~sumout ;
wire \add_sub_cella[9]~sumout ;
wire \add_sub_cella[10]~sumout ;


dffeas dffe18(
	.clk(clock),
	.d(\add_sub_cella[17]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe181),
	.prn(vcc));
defparam dffe18.is_wysiwyg = "true";
defparam dffe18.power_up = "low";

dffeas dffe17(
	.clk(clock),
	.d(\add_sub_cella[16]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe171),
	.prn(vcc));
defparam dffe17.is_wysiwyg = "true";
defparam dffe17.power_up = "low";

dffeas dffe16(
	.clk(clock),
	.d(\add_sub_cella[15]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe161),
	.prn(vcc));
defparam dffe16.is_wysiwyg = "true";
defparam dffe16.power_up = "low";

dffeas dffe15(
	.clk(clock),
	.d(\add_sub_cella[14]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe151),
	.prn(vcc));
defparam dffe15.is_wysiwyg = "true";
defparam dffe15.power_up = "low";

dffeas dffe14(
	.clk(clock),
	.d(\add_sub_cella[13]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe141),
	.prn(vcc));
defparam dffe14.is_wysiwyg = "true";
defparam dffe14.power_up = "low";

dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

dffeas dffe13(
	.clk(clock),
	.d(\add_sub_cella[12]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe131),
	.prn(vcc));
defparam dffe13.is_wysiwyg = "true";
defparam dffe13.power_up = "low";

dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe19),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

arriav_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_1),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_2),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_3),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_4),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_5),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_6),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(\add_sub_cella[11]~COUT ),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[12] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[11]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[12]~sumout ),
	.cout(\add_sub_cella[12]~COUT ),
	.shareout());
defparam \add_sub_cella[12] .extended_lut = "off";
defparam \add_sub_cella[12] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[12] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[13] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[12]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[13]~sumout ),
	.cout(\add_sub_cella[13]~COUT ),
	.shareout());
defparam \add_sub_cella[13] .extended_lut = "off";
defparam \add_sub_cella[13] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[13] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[14] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[13]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[14]~sumout ),
	.cout(\add_sub_cella[14]~COUT ),
	.shareout());
defparam \add_sub_cella[14] .extended_lut = "off";
defparam \add_sub_cella[14] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[14] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[15] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[14]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[15]~sumout ),
	.cout(\add_sub_cella[15]~COUT ),
	.shareout());
defparam \add_sub_cella[15] .extended_lut = "off";
defparam \add_sub_cella[15] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[15] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[16] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_16),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[15]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[16]~sumout ),
	.cout(\add_sub_cella[16]~COUT ),
	.shareout());
defparam \add_sub_cella[16] .extended_lut = "off";
defparam \add_sub_cella[16] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[16] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[17] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_17),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[16]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[17]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[17] .extended_lut = "off";
defparam \add_sub_cella[17] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[17] .shared_arith = "off";

endmodule

module nco_test_cordic_sxor_1p_lpm_8 (
	sin_o_0,
	dffe18,
	dffe17,
	dffe16,
	dffe161,
	dffe181,
	pipeline_dffe_17,
	dffe15,
	dffe13,
	dffe14,
	pipeline_dffe_16,
	dffe171,
	pipeline_dffe_15,
	dffe1,
	dffe162,
	dffe2,
	dffe3,
	dffe4,
	dffe5,
	dffe6,
	dffe7,
	dffe8,
	dffe9,
	dffe10,
	dffe11,
	dffe12,
	pipeline_dffe_14,
	dffe151,
	pipeline_dffe_13,
	dffe141,
	dffe121,
	dffe131,
	pipeline_dffe_12,
	pipeline_dffe_11,
	dffe19,
	dffe21,
	dffe31,
	dffe41,
	dffe51,
	dffe61,
	dffe71,
	dffe81,
	dffe91,
	dffe101,
	dffe111,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	sin_o_0;
output 	dffe18;
output 	dffe17;
input 	dffe16;
output 	dffe161;
input 	dffe181;
input 	pipeline_dffe_17;
output 	dffe15;
output 	dffe13;
output 	dffe14;
input 	pipeline_dffe_16;
input 	dffe171;
input 	pipeline_dffe_15;
output 	dffe1;
input 	dffe162;
output 	dffe2;
output 	dffe3;
output 	dffe4;
output 	dffe5;
output 	dffe6;
output 	dffe7;
output 	dffe8;
output 	dffe9;
output 	dffe10;
output 	dffe11;
output 	dffe12;
input 	pipeline_dffe_14;
input 	dffe151;
input 	pipeline_dffe_13;
input 	dffe141;
input 	dffe121;
input 	dffe131;
input 	pipeline_dffe_12;
input 	pipeline_dffe_11;
input 	dffe19;
input 	dffe21;
input 	dffe31;
input 	dffe41;
input 	dffe51;
input 	dffe61;
input 	dffe71;
input 	dffe81;
input 	dffe91;
input 	dffe101;
input 	dffe111;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[17]~q ;
wire \xordvalue[10]~q ;
wire \Add0~1_sumout ;
wire \a[16]~q ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \a[15]~q ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \a[14]~q ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \a[13]~q ;
wire \a[12]~q ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \a[11]~q ;
wire \a[0]~q ;
wire \xordvalue[0]~q ;
wire \a[1]~q ;
wire \xordvalue[1]~q ;
wire \a[2]~q ;
wire \xordvalue[2]~q ;
wire \a[3]~q ;
wire \xordvalue[3]~q ;
wire \a[4]~q ;
wire \xordvalue[4]~q ;
wire \a[5]~q ;
wire \xordvalue[5]~q ;
wire \a[6]~q ;
wire \a[7]~q ;
wire \a[8]~q ;
wire \a[9]~q ;
wire \a[10]~q ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~51 ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~55 ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~59 ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~63 ;
wire \Add0~65_sumout ;
wire \Add0~66 ;
wire \Add0~67 ;
wire \Add0~69_sumout ;
wire \Add0~70 ;
wire \Add0~71 ;
wire \xordvalue~0_combout ;
wire \xordvalue~1_combout ;
wire \xordvalue~2_combout ;
wire \xordvalue~3_combout ;
wire \xordvalue~4_combout ;
wire \xordvalue~5_combout ;
wire \xordvalue~6_combout ;


nco_test_lpm_add_sub_27 u0(
	.a_17(\a[17]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.a_16(\a[16]~q ),
	.a_15(\a[15]~q ),
	.a_14(\a[14]~q ),
	.a_13(\a[13]~q ),
	.a_12(\a[12]~q ),
	.a_11(\a[11]~q ),
	.a_0(\a[0]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_1(\a[1]~q ),
	.xordvalue_1(\xordvalue[1]~q ),
	.a_2(\a[2]~q ),
	.xordvalue_2(\xordvalue[2]~q ),
	.a_3(\a[3]~q ),
	.xordvalue_3(\xordvalue[3]~q ),
	.a_4(\a[4]~q ),
	.xordvalue_4(\xordvalue[4]~q ),
	.a_5(\a[5]~q ),
	.xordvalue_5(\xordvalue[5]~q ),
	.a_6(\a[6]~q ),
	.a_7(\a[7]~q ),
	.a_8(\a[8]~q ),
	.a_9(\a[9]~q ),
	.a_10(\a[10]~q ),
	.dffe18(dffe18),
	.dffe17(dffe17),
	.dffe16(dffe161),
	.dffe15(dffe15),
	.dffe13(dffe13),
	.dffe14(dffe14),
	.dffe1(dffe1),
	.dffe2(dffe2),
	.dffe3(dffe3),
	.dffe4(dffe4),
	.dffe5(dffe5),
	.dffe6(dffe6),
	.dffe7(dffe7),
	.dffe8(dffe8),
	.dffe9(dffe9),
	.dffe10(dffe10),
	.dffe11(dffe11),
	.dffe12(dffe12),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[17] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[17]~q ),
	.prn(vcc));
defparam \a[17] .is_wysiwyg = "true";
defparam \a[17] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe181),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "on";

dffeas \a[16] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[16]~q ),
	.prn(vcc));
defparam \a[16] .is_wysiwyg = "true";
defparam \a[16] .power_up = "low";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe171),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~5 .shared_arith = "on";

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe162),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~9 .shared_arith = "on";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~13 .shared_arith = "on";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~17 .shared_arith = "on";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "on";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \xordvalue[1] (
	.clk(clk),
	.d(\xordvalue~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[1]~q ),
	.prn(vcc));
defparam \xordvalue[1] .is_wysiwyg = "true";
defparam \xordvalue[1] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \xordvalue[2] (
	.clk(clk),
	.d(\xordvalue~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[2]~q ),
	.prn(vcc));
defparam \xordvalue[2] .is_wysiwyg = "true";
defparam \xordvalue[2] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \xordvalue[3] (
	.clk(clk),
	.d(\xordvalue~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[3]~q ),
	.prn(vcc));
defparam \xordvalue[3] .is_wysiwyg = "true";
defparam \xordvalue[3] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \xordvalue[4] (
	.clk(clk),
	.d(\xordvalue~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[4]~q ),
	.prn(vcc));
defparam \xordvalue[4] .is_wysiwyg = "true";
defparam \xordvalue[4] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \xordvalue[5] (
	.clk(clk),
	.d(\xordvalue~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[5]~q ),
	.prn(vcc));
defparam \xordvalue[5] .is_wysiwyg = "true";
defparam \xordvalue[5] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~70 ),
	.sharein(\Add0~71 ),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~25 .shared_arith = "on";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!dffe19),
	.datad(!dffe16),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add0~29 .shared_arith = "on";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~33 .shared_arith = "on";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~37 .shared_arith = "on";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~41 .shared_arith = "on";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout(\Add0~47 ));
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~45 .shared_arith = "on";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(\Add0~47 ),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout(\Add0~51 ));
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~49 .shared_arith = "on";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(\Add0~51 ),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout(\Add0~55 ));
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~53 .shared_arith = "on";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(\Add0~55 ),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout(\Add0~59 ));
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~57 .shared_arith = "on";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(\Add0~59 ),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout(\Add0~63 ));
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~61 .shared_arith = "on";

arriav_lcell_comb \Add0~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(\Add0~63 ),
	.combout(),
	.sumout(\Add0~65_sumout ),
	.cout(\Add0~66 ),
	.shareout(\Add0~67 ));
defparam \Add0~65 .extended_lut = "off";
defparam \Add0~65 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~65 .shared_arith = "on";

arriav_lcell_comb \Add0~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~66 ),
	.sharein(\Add0~67 ),
	.combout(),
	.sumout(\Add0~69_sumout ),
	.cout(\Add0~70 ),
	.shareout(\Add0~71 ));
defparam \Add0~69 .extended_lut = "off";
defparam \Add0~69 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~69 .shared_arith = "on";

arriav_lcell_comb \xordvalue~0 (
	.dataa(!pipeline_dffe_17),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

arriav_lcell_comb \xordvalue~1 (
	.dataa(!pipeline_dffe_11),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~1 .extended_lut = "off";
defparam \xordvalue~1 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~1 .shared_arith = "off";

arriav_lcell_comb \xordvalue~2 (
	.dataa(!pipeline_dffe_12),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~2 .extended_lut = "off";
defparam \xordvalue~2 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~2 .shared_arith = "off";

arriav_lcell_comb \xordvalue~3 (
	.dataa(!pipeline_dffe_13),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~3 .extended_lut = "off";
defparam \xordvalue~3 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~3 .shared_arith = "off";

arriav_lcell_comb \xordvalue~4 (
	.dataa(!pipeline_dffe_14),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~4 .extended_lut = "off";
defparam \xordvalue~4 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~4 .shared_arith = "off";

arriav_lcell_comb \xordvalue~5 (
	.dataa(!pipeline_dffe_15),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~5 .extended_lut = "off";
defparam \xordvalue~5 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~5 .shared_arith = "off";

arriav_lcell_comb \xordvalue~6 (
	.dataa(!pipeline_dffe_16),
	.datab(!dffe16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~6 .extended_lut = "off";
defparam \xordvalue~6 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~6 .shared_arith = "off";

endmodule

module nco_test_lpm_add_sub_27 (
	a_17,
	xordvalue_10,
	a_16,
	a_15,
	a_14,
	a_13,
	a_12,
	a_11,
	a_0,
	xordvalue_0,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	a_4,
	xordvalue_4,
	a_5,
	xordvalue_5,
	a_6,
	a_7,
	a_8,
	a_9,
	a_10,
	dffe18,
	dffe17,
	dffe16,
	dffe15,
	dffe13,
	dffe14,
	dffe1,
	dffe2,
	dffe3,
	dffe4,
	dffe5,
	dffe6,
	dffe7,
	dffe8,
	dffe9,
	dffe10,
	dffe11,
	dffe12,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_10;
input 	a_16;
input 	a_15;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_0;
input 	xordvalue_0;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
input 	a_4;
input 	xordvalue_4;
input 	a_5;
input 	xordvalue_5;
input 	a_6;
input 	a_7;
input 	a_8;
input 	a_9;
input 	a_10;
output 	dffe18;
output 	dffe17;
output 	dffe16;
output 	dffe15;
output 	dffe13;
output 	dffe14;
output 	dffe1;
output 	dffe2;
output 	dffe3;
output 	dffe4;
output 	dffe5;
output 	dffe6;
output 	dffe7;
output 	dffe8;
output 	dffe9;
output 	dffe10;
output 	dffe11;
output 	dffe12;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_add_sub_jdg_8 auto_generated(
	.a_17(a_17),
	.xordvalue_10(xordvalue_10),
	.a_16(a_16),
	.a_15(a_15),
	.a_14(a_14),
	.a_13(a_13),
	.a_12(a_12),
	.a_11(a_11),
	.a_0(a_0),
	.xordvalue_0(xordvalue_0),
	.a_1(a_1),
	.xordvalue_1(xordvalue_1),
	.a_2(a_2),
	.xordvalue_2(xordvalue_2),
	.a_3(a_3),
	.xordvalue_3(xordvalue_3),
	.a_4(a_4),
	.xordvalue_4(xordvalue_4),
	.a_5(a_5),
	.xordvalue_5(xordvalue_5),
	.a_6(a_6),
	.a_7(a_7),
	.a_8(a_8),
	.a_9(a_9),
	.a_10(a_10),
	.dffe181(dffe18),
	.dffe171(dffe17),
	.dffe161(dffe16),
	.dffe151(dffe15),
	.dffe131(dffe13),
	.dffe141(dffe14),
	.dffe19(dffe1),
	.dffe21(dffe2),
	.dffe31(dffe3),
	.dffe41(dffe4),
	.dffe51(dffe5),
	.dffe61(dffe6),
	.dffe71(dffe7),
	.dffe81(dffe8),
	.dffe91(dffe9),
	.dffe101(dffe10),
	.dffe111(dffe11),
	.dffe121(dffe12),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module nco_test_add_sub_jdg_8 (
	a_17,
	xordvalue_10,
	a_16,
	a_15,
	a_14,
	a_13,
	a_12,
	a_11,
	a_0,
	xordvalue_0,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	a_4,
	xordvalue_4,
	a_5,
	xordvalue_5,
	a_6,
	a_7,
	a_8,
	a_9,
	a_10,
	dffe181,
	dffe171,
	dffe161,
	dffe151,
	dffe131,
	dffe141,
	dffe19,
	dffe21,
	dffe31,
	dffe41,
	dffe51,
	dffe61,
	dffe71,
	dffe81,
	dffe91,
	dffe101,
	dffe111,
	dffe121,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_10;
input 	a_16;
input 	a_15;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_0;
input 	xordvalue_0;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
input 	a_4;
input 	xordvalue_4;
input 	a_5;
input 	xordvalue_5;
input 	a_6;
input 	a_7;
input 	a_8;
input 	a_9;
input 	a_10;
output 	dffe181;
output 	dffe171;
output 	dffe161;
output 	dffe151;
output 	dffe131;
output 	dffe141;
output 	dffe19;
output 	dffe21;
output 	dffe31;
output 	dffe41;
output 	dffe51;
output 	dffe61;
output 	dffe71;
output 	dffe81;
output 	dffe91;
output 	dffe101;
output 	dffe111;
output 	dffe121;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~COUT ;
wire \add_sub_cella[12]~COUT ;
wire \add_sub_cella[13]~COUT ;
wire \add_sub_cella[14]~COUT ;
wire \add_sub_cella[15]~COUT ;
wire \add_sub_cella[16]~COUT ;
wire \add_sub_cella[17]~sumout ;
wire \add_sub_cella[16]~sumout ;
wire \add_sub_cella[15]~sumout ;
wire \add_sub_cella[14]~sumout ;
wire \add_sub_cella[12]~sumout ;
wire \add_sub_cella[13]~sumout ;
wire \add_sub_cella[0]~sumout ;
wire \add_sub_cella[1]~sumout ;
wire \add_sub_cella[2]~sumout ;
wire \add_sub_cella[3]~sumout ;
wire \add_sub_cella[4]~sumout ;
wire \add_sub_cella[5]~sumout ;
wire \add_sub_cella[6]~sumout ;
wire \add_sub_cella[7]~sumout ;
wire \add_sub_cella[8]~sumout ;
wire \add_sub_cella[9]~sumout ;
wire \add_sub_cella[10]~sumout ;
wire \add_sub_cella[11]~sumout ;


dffeas dffe18(
	.clk(clock),
	.d(\add_sub_cella[17]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe181),
	.prn(vcc));
defparam dffe18.is_wysiwyg = "true";
defparam dffe18.power_up = "low";

dffeas dffe17(
	.clk(clock),
	.d(\add_sub_cella[16]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe171),
	.prn(vcc));
defparam dffe17.is_wysiwyg = "true";
defparam dffe17.power_up = "low";

dffeas dffe16(
	.clk(clock),
	.d(\add_sub_cella[15]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe161),
	.prn(vcc));
defparam dffe16.is_wysiwyg = "true";
defparam dffe16.power_up = "low";

dffeas dffe15(
	.clk(clock),
	.d(\add_sub_cella[14]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe151),
	.prn(vcc));
defparam dffe15.is_wysiwyg = "true";
defparam dffe15.power_up = "low";

dffeas dffe13(
	.clk(clock),
	.d(\add_sub_cella[12]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe131),
	.prn(vcc));
defparam dffe13.is_wysiwyg = "true";
defparam dffe13.power_up = "low";

dffeas dffe14(
	.clk(clock),
	.d(\add_sub_cella[13]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe141),
	.prn(vcc));
defparam dffe14.is_wysiwyg = "true";
defparam dffe14.power_up = "low";

dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe19),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

arriav_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_1),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_2),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_3),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_4),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_5),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(\add_sub_cella[11]~COUT ),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[12] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[11]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[12]~sumout ),
	.cout(\add_sub_cella[12]~COUT ),
	.shareout());
defparam \add_sub_cella[12] .extended_lut = "off";
defparam \add_sub_cella[12] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[12] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[13] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[12]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[13]~sumout ),
	.cout(\add_sub_cella[13]~COUT ),
	.shareout());
defparam \add_sub_cella[13] .extended_lut = "off";
defparam \add_sub_cella[13] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[13] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[14] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[13]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[14]~sumout ),
	.cout(\add_sub_cella[14]~COUT ),
	.shareout());
defparam \add_sub_cella[14] .extended_lut = "off";
defparam \add_sub_cella[14] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[14] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[15] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[14]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[15]~sumout ),
	.cout(\add_sub_cella[15]~COUT ),
	.shareout());
defparam \add_sub_cella[15] .extended_lut = "off";
defparam \add_sub_cella[15] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[15] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[16] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_16),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[15]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[16]~sumout ),
	.cout(\add_sub_cella[16]~COUT ),
	.shareout());
defparam \add_sub_cella[16] .extended_lut = "off";
defparam \add_sub_cella[16] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[16] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[17] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_17),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[16]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[17]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[17] .extended_lut = "off";
defparam \add_sub_cella[17] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[17] .shared_arith = "off";

endmodule

module nco_test_cordic_sxor_1p_lpm_9 (
	sin_o_0,
	dffe18,
	dffe17,
	dffe16,
	pipeline_dffe_17,
	dffe161,
	dffe181,
	dffe14,
	dffe15,
	dffe171,
	dffe1,
	pipeline_dffe_16,
	dffe2,
	dffe3,
	dffe4,
	dffe5,
	dffe6,
	dffe7,
	dffe8,
	dffe9,
	dffe10,
	dffe11,
	dffe12,
	dffe13,
	dffe162,
	pipeline_dffe_15,
	dffe151,
	pipeline_dffe_14,
	dffe131,
	dffe141,
	pipeline_dffe_12,
	pipeline_dffe_13,
	dffe19,
	dffe21,
	dffe31,
	dffe41,
	dffe51,
	dffe61,
	dffe71,
	dffe81,
	dffe91,
	dffe101,
	dffe111,
	dffe121,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	sin_o_0;
output 	dffe18;
output 	dffe17;
input 	dffe16;
input 	pipeline_dffe_17;
output 	dffe161;
input 	dffe181;
output 	dffe14;
output 	dffe15;
input 	dffe171;
output 	dffe1;
input 	pipeline_dffe_16;
output 	dffe2;
output 	dffe3;
output 	dffe4;
output 	dffe5;
output 	dffe6;
output 	dffe7;
output 	dffe8;
output 	dffe9;
output 	dffe10;
output 	dffe11;
output 	dffe12;
output 	dffe13;
input 	dffe162;
input 	pipeline_dffe_15;
input 	dffe151;
input 	pipeline_dffe_14;
input 	dffe131;
input 	dffe141;
input 	pipeline_dffe_12;
input 	pipeline_dffe_13;
input 	dffe19;
input 	dffe21;
input 	dffe31;
input 	dffe41;
input 	dffe51;
input 	dffe61;
input 	dffe71;
input 	dffe81;
input 	dffe91;
input 	dffe101;
input 	dffe111;
input 	dffe121;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[17]~q ;
wire \xordvalue[10]~q ;
wire \Add0~1_sumout ;
wire \a[16]~q ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \a[15]~q ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \a[14]~q ;
wire \a[13]~q ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \a[12]~q ;
wire \a[0]~q ;
wire \xordvalue[0]~q ;
wire \a[1]~q ;
wire \xordvalue[1]~q ;
wire \a[2]~q ;
wire \xordvalue[2]~q ;
wire \a[3]~q ;
wire \xordvalue[3]~q ;
wire \a[4]~q ;
wire \xordvalue[4]~q ;
wire \a[5]~q ;
wire \a[6]~q ;
wire \a[7]~q ;
wire \a[8]~q ;
wire \a[9]~q ;
wire \a[10]~q ;
wire \a[11]~q ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~51 ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~55 ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~59 ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~63 ;
wire \Add0~65_sumout ;
wire \Add0~66 ;
wire \Add0~67 ;
wire \Add0~69_sumout ;
wire \Add0~70 ;
wire \Add0~71 ;
wire \xordvalue~0_combout ;
wire \xordvalue~1_combout ;
wire \xordvalue~2_combout ;
wire \xordvalue~3_combout ;
wire \xordvalue~4_combout ;
wire \xordvalue~5_combout ;


nco_test_lpm_add_sub_28 u0(
	.a_17(\a[17]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.a_16(\a[16]~q ),
	.a_15(\a[15]~q ),
	.a_14(\a[14]~q ),
	.a_13(\a[13]~q ),
	.a_12(\a[12]~q ),
	.a_0(\a[0]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_1(\a[1]~q ),
	.xordvalue_1(\xordvalue[1]~q ),
	.a_2(\a[2]~q ),
	.xordvalue_2(\xordvalue[2]~q ),
	.a_3(\a[3]~q ),
	.xordvalue_3(\xordvalue[3]~q ),
	.a_4(\a[4]~q ),
	.xordvalue_4(\xordvalue[4]~q ),
	.a_5(\a[5]~q ),
	.a_6(\a[6]~q ),
	.a_7(\a[7]~q ),
	.a_8(\a[8]~q ),
	.a_9(\a[9]~q ),
	.a_10(\a[10]~q ),
	.a_11(\a[11]~q ),
	.dffe18(dffe18),
	.dffe17(dffe17),
	.dffe16(dffe161),
	.dffe14(dffe14),
	.dffe15(dffe15),
	.dffe1(dffe1),
	.dffe2(dffe2),
	.dffe3(dffe3),
	.dffe4(dffe4),
	.dffe5(dffe5),
	.dffe6(dffe6),
	.dffe7(dffe7),
	.dffe8(dffe8),
	.dffe9(dffe9),
	.dffe10(dffe10),
	.dffe11(dffe11),
	.dffe12(dffe12),
	.dffe13(dffe13),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[17] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[17]~q ),
	.prn(vcc));
defparam \a[17] .is_wysiwyg = "true";
defparam \a[17] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe181),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "on";

dffeas \a[16] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[16]~q ),
	.prn(vcc));
defparam \a[16] .is_wysiwyg = "true";
defparam \a[16] .power_up = "low";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe171),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~5 .shared_arith = "on";

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe162),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~9 .shared_arith = "on";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~13 .shared_arith = "on";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~17 .shared_arith = "on";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \xordvalue[1] (
	.clk(clk),
	.d(\xordvalue~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[1]~q ),
	.prn(vcc));
defparam \xordvalue[1] .is_wysiwyg = "true";
defparam \xordvalue[1] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \xordvalue[2] (
	.clk(clk),
	.d(\xordvalue~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[2]~q ),
	.prn(vcc));
defparam \xordvalue[2] .is_wysiwyg = "true";
defparam \xordvalue[2] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \xordvalue[3] (
	.clk(clk),
	.d(\xordvalue~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[3]~q ),
	.prn(vcc));
defparam \xordvalue[3] .is_wysiwyg = "true";
defparam \xordvalue[3] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \xordvalue[4] (
	.clk(clk),
	.d(\xordvalue~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[4]~q ),
	.prn(vcc));
defparam \xordvalue[4] .is_wysiwyg = "true";
defparam \xordvalue[4] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~70 ),
	.sharein(\Add0~71 ),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "on";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!dffe19),
	.datad(!dffe16),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add0~25 .shared_arith = "on";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~29 .shared_arith = "on";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~33 .shared_arith = "on";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~37 .shared_arith = "on";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~41 .shared_arith = "on";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout(\Add0~47 ));
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~45 .shared_arith = "on";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(\Add0~47 ),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout(\Add0~51 ));
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~49 .shared_arith = "on";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(\Add0~51 ),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout(\Add0~55 ));
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~53 .shared_arith = "on";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(\Add0~55 ),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout(\Add0~59 ));
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~57 .shared_arith = "on";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(\Add0~59 ),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout(\Add0~63 ));
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~61 .shared_arith = "on";

arriav_lcell_comb \Add0~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(\Add0~63 ),
	.combout(),
	.sumout(\Add0~65_sumout ),
	.cout(\Add0~66 ),
	.shareout(\Add0~67 ));
defparam \Add0~65 .extended_lut = "off";
defparam \Add0~65 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~65 .shared_arith = "on";

arriav_lcell_comb \Add0~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~66 ),
	.sharein(\Add0~67 ),
	.combout(),
	.sumout(\Add0~69_sumout ),
	.cout(\Add0~70 ),
	.shareout(\Add0~71 ));
defparam \Add0~69 .extended_lut = "off";
defparam \Add0~69 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~69 .shared_arith = "on";

arriav_lcell_comb \xordvalue~0 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_17),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

arriav_lcell_comb \xordvalue~1 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_12),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~1 .extended_lut = "off";
defparam \xordvalue~1 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~1 .shared_arith = "off";

arriav_lcell_comb \xordvalue~2 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_13),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~2 .extended_lut = "off";
defparam \xordvalue~2 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~2 .shared_arith = "off";

arriav_lcell_comb \xordvalue~3 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_14),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~3 .extended_lut = "off";
defparam \xordvalue~3 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~3 .shared_arith = "off";

arriav_lcell_comb \xordvalue~4 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_15),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~4 .extended_lut = "off";
defparam \xordvalue~4 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~4 .shared_arith = "off";

arriav_lcell_comb \xordvalue~5 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~5 .extended_lut = "off";
defparam \xordvalue~5 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~5 .shared_arith = "off";

endmodule

module nco_test_lpm_add_sub_28 (
	a_17,
	xordvalue_10,
	a_16,
	a_15,
	a_14,
	a_13,
	a_12,
	a_0,
	xordvalue_0,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	a_4,
	xordvalue_4,
	a_5,
	a_6,
	a_7,
	a_8,
	a_9,
	a_10,
	a_11,
	dffe18,
	dffe17,
	dffe16,
	dffe14,
	dffe15,
	dffe1,
	dffe2,
	dffe3,
	dffe4,
	dffe5,
	dffe6,
	dffe7,
	dffe8,
	dffe9,
	dffe10,
	dffe11,
	dffe12,
	dffe13,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_10;
input 	a_16;
input 	a_15;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_0;
input 	xordvalue_0;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
input 	a_4;
input 	xordvalue_4;
input 	a_5;
input 	a_6;
input 	a_7;
input 	a_8;
input 	a_9;
input 	a_10;
input 	a_11;
output 	dffe18;
output 	dffe17;
output 	dffe16;
output 	dffe14;
output 	dffe15;
output 	dffe1;
output 	dffe2;
output 	dffe3;
output 	dffe4;
output 	dffe5;
output 	dffe6;
output 	dffe7;
output 	dffe8;
output 	dffe9;
output 	dffe10;
output 	dffe11;
output 	dffe12;
output 	dffe13;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_add_sub_jdg_9 auto_generated(
	.a_17(a_17),
	.xordvalue_10(xordvalue_10),
	.a_16(a_16),
	.a_15(a_15),
	.a_14(a_14),
	.a_13(a_13),
	.a_12(a_12),
	.a_0(a_0),
	.xordvalue_0(xordvalue_0),
	.a_1(a_1),
	.xordvalue_1(xordvalue_1),
	.a_2(a_2),
	.xordvalue_2(xordvalue_2),
	.a_3(a_3),
	.xordvalue_3(xordvalue_3),
	.a_4(a_4),
	.xordvalue_4(xordvalue_4),
	.a_5(a_5),
	.a_6(a_6),
	.a_7(a_7),
	.a_8(a_8),
	.a_9(a_9),
	.a_10(a_10),
	.a_11(a_11),
	.dffe181(dffe18),
	.dffe171(dffe17),
	.dffe161(dffe16),
	.dffe141(dffe14),
	.dffe151(dffe15),
	.dffe19(dffe1),
	.dffe21(dffe2),
	.dffe31(dffe3),
	.dffe41(dffe4),
	.dffe51(dffe5),
	.dffe61(dffe6),
	.dffe71(dffe7),
	.dffe81(dffe8),
	.dffe91(dffe9),
	.dffe101(dffe10),
	.dffe111(dffe11),
	.dffe121(dffe12),
	.dffe131(dffe13),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module nco_test_add_sub_jdg_9 (
	a_17,
	xordvalue_10,
	a_16,
	a_15,
	a_14,
	a_13,
	a_12,
	a_0,
	xordvalue_0,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	a_4,
	xordvalue_4,
	a_5,
	a_6,
	a_7,
	a_8,
	a_9,
	a_10,
	a_11,
	dffe181,
	dffe171,
	dffe161,
	dffe141,
	dffe151,
	dffe19,
	dffe21,
	dffe31,
	dffe41,
	dffe51,
	dffe61,
	dffe71,
	dffe81,
	dffe91,
	dffe101,
	dffe111,
	dffe121,
	dffe131,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_10;
input 	a_16;
input 	a_15;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_0;
input 	xordvalue_0;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
input 	a_4;
input 	xordvalue_4;
input 	a_5;
input 	a_6;
input 	a_7;
input 	a_8;
input 	a_9;
input 	a_10;
input 	a_11;
output 	dffe181;
output 	dffe171;
output 	dffe161;
output 	dffe141;
output 	dffe151;
output 	dffe19;
output 	dffe21;
output 	dffe31;
output 	dffe41;
output 	dffe51;
output 	dffe61;
output 	dffe71;
output 	dffe81;
output 	dffe91;
output 	dffe101;
output 	dffe111;
output 	dffe121;
output 	dffe131;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~COUT ;
wire \add_sub_cella[12]~COUT ;
wire \add_sub_cella[13]~COUT ;
wire \add_sub_cella[14]~COUT ;
wire \add_sub_cella[15]~COUT ;
wire \add_sub_cella[16]~COUT ;
wire \add_sub_cella[17]~sumout ;
wire \add_sub_cella[16]~sumout ;
wire \add_sub_cella[15]~sumout ;
wire \add_sub_cella[13]~sumout ;
wire \add_sub_cella[14]~sumout ;
wire \add_sub_cella[0]~sumout ;
wire \add_sub_cella[1]~sumout ;
wire \add_sub_cella[2]~sumout ;
wire \add_sub_cella[3]~sumout ;
wire \add_sub_cella[4]~sumout ;
wire \add_sub_cella[5]~sumout ;
wire \add_sub_cella[6]~sumout ;
wire \add_sub_cella[7]~sumout ;
wire \add_sub_cella[8]~sumout ;
wire \add_sub_cella[9]~sumout ;
wire \add_sub_cella[10]~sumout ;
wire \add_sub_cella[11]~sumout ;
wire \add_sub_cella[12]~sumout ;


dffeas dffe18(
	.clk(clock),
	.d(\add_sub_cella[17]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe181),
	.prn(vcc));
defparam dffe18.is_wysiwyg = "true";
defparam dffe18.power_up = "low";

dffeas dffe17(
	.clk(clock),
	.d(\add_sub_cella[16]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe171),
	.prn(vcc));
defparam dffe17.is_wysiwyg = "true";
defparam dffe17.power_up = "low";

dffeas dffe16(
	.clk(clock),
	.d(\add_sub_cella[15]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe161),
	.prn(vcc));
defparam dffe16.is_wysiwyg = "true";
defparam dffe16.power_up = "low";

dffeas dffe14(
	.clk(clock),
	.d(\add_sub_cella[13]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe141),
	.prn(vcc));
defparam dffe14.is_wysiwyg = "true";
defparam dffe14.power_up = "low";

dffeas dffe15(
	.clk(clock),
	.d(\add_sub_cella[14]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe151),
	.prn(vcc));
defparam dffe15.is_wysiwyg = "true";
defparam dffe15.power_up = "low";

dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe19),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

dffeas dffe13(
	.clk(clock),
	.d(\add_sub_cella[12]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe131),
	.prn(vcc));
defparam dffe13.is_wysiwyg = "true";
defparam dffe13.power_up = "low";

arriav_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_1),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_2),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_3),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_4),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(\add_sub_cella[11]~COUT ),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[12] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[11]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[12]~sumout ),
	.cout(\add_sub_cella[12]~COUT ),
	.shareout());
defparam \add_sub_cella[12] .extended_lut = "off";
defparam \add_sub_cella[12] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[12] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[13] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[12]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[13]~sumout ),
	.cout(\add_sub_cella[13]~COUT ),
	.shareout());
defparam \add_sub_cella[13] .extended_lut = "off";
defparam \add_sub_cella[13] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[13] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[14] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[13]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[14]~sumout ),
	.cout(\add_sub_cella[14]~COUT ),
	.shareout());
defparam \add_sub_cella[14] .extended_lut = "off";
defparam \add_sub_cella[14] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[14] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[15] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[14]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[15]~sumout ),
	.cout(\add_sub_cella[15]~COUT ),
	.shareout());
defparam \add_sub_cella[15] .extended_lut = "off";
defparam \add_sub_cella[15] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[15] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[16] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_16),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[15]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[16]~sumout ),
	.cout(\add_sub_cella[16]~COUT ),
	.shareout());
defparam \add_sub_cella[16] .extended_lut = "off";
defparam \add_sub_cella[16] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[16] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[17] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_17),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[16]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[17]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[17] .extended_lut = "off";
defparam \add_sub_cella[17] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[17] .shared_arith = "off";

endmodule

module nco_test_cordic_sxor_1p_lpm_10 (
	a_0,
	xordvalue_11,
	cor1x_10,
	sin_o_0,
	dffe18,
	dffe17,
	dffe16,
	xordvalue,
	dffe161,
	dffe15,
	dffe14,
	dffe13,
	dffe12,
	dffe11,
	dffe10,
	dffe9,
	dffe8,
	dffe7,
	dffe6,
	dffe5,
	dffe3,
	dffe4,
	dffe1,
	dffe2,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_0;
input 	xordvalue_11;
input 	cor1x_10;
input 	sin_o_0;
output 	dffe18;
output 	dffe17;
input 	dffe16;
input 	xordvalue;
output 	dffe161;
output 	dffe15;
output 	dffe14;
output 	dffe13;
output 	dffe12;
output 	dffe11;
output 	dffe10;
output 	dffe9;
output 	dffe8;
output 	dffe7;
output 	dffe6;
output 	dffe5;
output 	dffe3;
output 	dffe4;
output 	dffe1;
output 	dffe2;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[17]~q ;
wire \a[16]~q ;
wire \a[15]~q ;
wire \a[14]~q ;
wire \a[13]~q ;
wire \a[12]~q ;
wire \a[11]~q ;
wire \a[10]~q ;
wire \a[9]~q ;
wire \a[8]~q ;
wire \a[7]~q ;
wire \a[6]~q ;
wire \a[5]~q ;
wire \a[4]~q ;
wire \a[3]~q ;
wire \a[2]~q ;
wire \a[1]~q ;
wire \a[0]~q ;
wire \Add0~0_combout ;
wire \Add0~1_combout ;


nco_test_lpm_add_sub_33 u0(
	.a_0(a_0),
	.xordvalue_11(xordvalue_11),
	.a_17(\a[17]~q ),
	.a_16(\a[16]~q ),
	.a_15(\a[15]~q ),
	.a_14(\a[14]~q ),
	.a_13(\a[13]~q ),
	.a_12(\a[12]~q ),
	.a_11(\a[11]~q ),
	.a_10(\a[10]~q ),
	.a_9(\a[9]~q ),
	.a_8(\a[8]~q ),
	.a_7(\a[7]~q ),
	.a_6(\a[6]~q ),
	.a_5(\a[5]~q ),
	.a_4(\a[4]~q ),
	.a_3(\a[3]~q ),
	.a_2(\a[2]~q ),
	.a_1(\a[1]~q ),
	.a_01(\a[0]~q ),
	.dffe18(dffe18),
	.dffe17(dffe17),
	.dffe16(dffe161),
	.dffe15(dffe15),
	.dffe14(dffe14),
	.dffe13(dffe13),
	.dffe12(dffe12),
	.dffe11(dffe11),
	.dffe10(dffe10),
	.dffe9(dffe9),
	.dffe8(dffe8),
	.dffe7(dffe7),
	.dffe6(dffe6),
	.dffe5(dffe5),
	.dffe3(dffe3),
	.dffe4(dffe4),
	.dffe1(dffe1),
	.dffe2(dffe2),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[17] (
	.clk(clk),
	.d(\Add0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[17]~q ),
	.prn(vcc));
defparam \a[17] .is_wysiwyg = "true";
defparam \a[17] .power_up = "low";

dffeas \a[16] (
	.clk(clk),
	.d(\Add0~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[16]~q ),
	.prn(vcc));
defparam \a[16] .is_wysiwyg = "true";
defparam \a[16] .power_up = "low";

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(xordvalue),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(dffe16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(dffe16),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

arriav_lcell_comb \Add0~0 (
	.dataa(!dffe16),
	.datab(!cor1x_10),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~0 .extended_lut = "off";
defparam \Add0~0 .lut_mask = 64'hDDDDDDDDDDDDDDDD;
defparam \Add0~0 .shared_arith = "off";

arriav_lcell_comb \Add0~1 (
	.dataa(!dffe16),
	.datab(!cor1x_10),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\Add0~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h7777777777777777;
defparam \Add0~1 .shared_arith = "off";

endmodule

module nco_test_cordic_sxor_1p_lpm_11 (
	sin_o_0,
	dffe18,
	dffe17,
	dffe15,
	dffe16,
	dffe161,
	dffe181,
	pipeline_dffe_17,
	dffe1,
	dffe2,
	dffe3,
	dffe4,
	dffe5,
	dffe6,
	dffe7,
	dffe8,
	dffe9,
	dffe10,
	dffe11,
	dffe12,
	dffe13,
	dffe14,
	pipeline_dffe_16,
	dffe171,
	pipeline_dffe_15,
	dffe162,
	dffe141,
	dffe151,
	pipeline_dffe_14,
	pipeline_dffe_13,
	dffe19,
	dffe21,
	dffe31,
	dffe41,
	dffe51,
	dffe61,
	dffe71,
	dffe81,
	dffe91,
	dffe101,
	dffe111,
	dffe121,
	dffe131,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	sin_o_0;
output 	dffe18;
output 	dffe17;
output 	dffe15;
output 	dffe16;
input 	dffe161;
input 	dffe181;
input 	pipeline_dffe_17;
output 	dffe1;
output 	dffe2;
output 	dffe3;
output 	dffe4;
output 	dffe5;
output 	dffe6;
output 	dffe7;
output 	dffe8;
output 	dffe9;
output 	dffe10;
output 	dffe11;
output 	dffe12;
output 	dffe13;
output 	dffe14;
input 	pipeline_dffe_16;
input 	dffe171;
input 	pipeline_dffe_15;
input 	dffe162;
input 	dffe141;
input 	dffe151;
input 	pipeline_dffe_14;
input 	pipeline_dffe_13;
input 	dffe19;
input 	dffe21;
input 	dffe31;
input 	dffe41;
input 	dffe51;
input 	dffe61;
input 	dffe71;
input 	dffe81;
input 	dffe91;
input 	dffe101;
input 	dffe111;
input 	dffe121;
input 	dffe131;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[17]~q ;
wire \xordvalue[10]~q ;
wire \Add0~1_sumout ;
wire \a[16]~q ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \a[15]~q ;
wire \a[14]~q ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \a[13]~q ;
wire \a[0]~q ;
wire \xordvalue[0]~q ;
wire \a[1]~q ;
wire \xordvalue[1]~q ;
wire \a[2]~q ;
wire \xordvalue[2]~q ;
wire \a[3]~q ;
wire \xordvalue[3]~q ;
wire \a[4]~q ;
wire \a[5]~q ;
wire \a[6]~q ;
wire \a[7]~q ;
wire \a[8]~q ;
wire \a[9]~q ;
wire \a[10]~q ;
wire \a[11]~q ;
wire \a[12]~q ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~51 ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~55 ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~59 ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~63 ;
wire \Add0~65_sumout ;
wire \Add0~66 ;
wire \Add0~67 ;
wire \Add0~69_sumout ;
wire \Add0~70 ;
wire \Add0~71 ;
wire \xordvalue~0_combout ;
wire \xordvalue~1_combout ;
wire \xordvalue~2_combout ;
wire \xordvalue~3_combout ;
wire \xordvalue~4_combout ;


nco_test_lpm_add_sub_29 u0(
	.a_17(\a[17]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.a_16(\a[16]~q ),
	.a_15(\a[15]~q ),
	.a_14(\a[14]~q ),
	.a_13(\a[13]~q ),
	.a_0(\a[0]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_1(\a[1]~q ),
	.xordvalue_1(\xordvalue[1]~q ),
	.a_2(\a[2]~q ),
	.xordvalue_2(\xordvalue[2]~q ),
	.a_3(\a[3]~q ),
	.xordvalue_3(\xordvalue[3]~q ),
	.a_4(\a[4]~q ),
	.a_5(\a[5]~q ),
	.a_6(\a[6]~q ),
	.a_7(\a[7]~q ),
	.a_8(\a[8]~q ),
	.a_9(\a[9]~q ),
	.a_10(\a[10]~q ),
	.a_11(\a[11]~q ),
	.a_12(\a[12]~q ),
	.dffe18(dffe18),
	.dffe17(dffe17),
	.dffe15(dffe15),
	.dffe16(dffe16),
	.dffe1(dffe1),
	.dffe2(dffe2),
	.dffe3(dffe3),
	.dffe4(dffe4),
	.dffe5(dffe5),
	.dffe6(dffe6),
	.dffe7(dffe7),
	.dffe8(dffe8),
	.dffe9(dffe9),
	.dffe10(dffe10),
	.dffe11(dffe11),
	.dffe12(dffe12),
	.dffe13(dffe13),
	.dffe14(dffe14),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[17] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[17]~q ),
	.prn(vcc));
defparam \a[17] .is_wysiwyg = "true";
defparam \a[17] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe181),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "on";

dffeas \a[16] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[16]~q ),
	.prn(vcc));
defparam \a[16] .is_wysiwyg = "true";
defparam \a[16] .power_up = "low";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe171),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~5 .shared_arith = "on";

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe162),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~9 .shared_arith = "on";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~13 .shared_arith = "on";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \xordvalue[1] (
	.clk(clk),
	.d(\xordvalue~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[1]~q ),
	.prn(vcc));
defparam \xordvalue[1] .is_wysiwyg = "true";
defparam \xordvalue[1] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \xordvalue[2] (
	.clk(clk),
	.d(\xordvalue~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[2]~q ),
	.prn(vcc));
defparam \xordvalue[2] .is_wysiwyg = "true";
defparam \xordvalue[2] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \xordvalue[3] (
	.clk(clk),
	.d(\xordvalue~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[3]~q ),
	.prn(vcc));
defparam \xordvalue[3] .is_wysiwyg = "true";
defparam \xordvalue[3] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~70 ),
	.sharein(\Add0~71 ),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~17 .shared_arith = "on";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!dffe19),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add0~21 .shared_arith = "on";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~25 .shared_arith = "on";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~29 .shared_arith = "on";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~33 .shared_arith = "on";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~37 .shared_arith = "on";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~41 .shared_arith = "on";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout(\Add0~47 ));
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~45 .shared_arith = "on";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(\Add0~47 ),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout(\Add0~51 ));
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~49 .shared_arith = "on";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(\Add0~51 ),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout(\Add0~55 ));
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~53 .shared_arith = "on";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(\Add0~55 ),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout(\Add0~59 ));
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~57 .shared_arith = "on";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(\Add0~59 ),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout(\Add0~63 ));
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~61 .shared_arith = "on";

arriav_lcell_comb \Add0~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(\Add0~63 ),
	.combout(),
	.sumout(\Add0~65_sumout ),
	.cout(\Add0~66 ),
	.shareout(\Add0~67 ));
defparam \Add0~65 .extended_lut = "off";
defparam \Add0~65 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~65 .shared_arith = "on";

arriav_lcell_comb \Add0~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~66 ),
	.sharein(\Add0~67 ),
	.combout(),
	.sumout(\Add0~69_sumout ),
	.cout(\Add0~70 ),
	.shareout(\Add0~71 ));
defparam \Add0~69 .extended_lut = "off";
defparam \Add0~69 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~69 .shared_arith = "on";

arriav_lcell_comb \xordvalue~0 (
	.dataa(!pipeline_dffe_17),
	.datab(!dffe161),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

arriav_lcell_comb \xordvalue~1 (
	.dataa(!pipeline_dffe_13),
	.datab(!dffe161),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~1 .extended_lut = "off";
defparam \xordvalue~1 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~1 .shared_arith = "off";

arriav_lcell_comb \xordvalue~2 (
	.dataa(!pipeline_dffe_14),
	.datab(!dffe161),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~2 .extended_lut = "off";
defparam \xordvalue~2 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~2 .shared_arith = "off";

arriav_lcell_comb \xordvalue~3 (
	.dataa(!pipeline_dffe_15),
	.datab(!dffe161),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~3 .extended_lut = "off";
defparam \xordvalue~3 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~3 .shared_arith = "off";

arriav_lcell_comb \xordvalue~4 (
	.dataa(!pipeline_dffe_16),
	.datab(!dffe161),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~4 .extended_lut = "off";
defparam \xordvalue~4 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~4 .shared_arith = "off";

endmodule

module nco_test_lpm_add_sub_29 (
	a_17,
	xordvalue_10,
	a_16,
	a_15,
	a_14,
	a_13,
	a_0,
	xordvalue_0,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	a_4,
	a_5,
	a_6,
	a_7,
	a_8,
	a_9,
	a_10,
	a_11,
	a_12,
	dffe18,
	dffe17,
	dffe15,
	dffe16,
	dffe1,
	dffe2,
	dffe3,
	dffe4,
	dffe5,
	dffe6,
	dffe7,
	dffe8,
	dffe9,
	dffe10,
	dffe11,
	dffe12,
	dffe13,
	dffe14,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_10;
input 	a_16;
input 	a_15;
input 	a_14;
input 	a_13;
input 	a_0;
input 	xordvalue_0;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
input 	a_4;
input 	a_5;
input 	a_6;
input 	a_7;
input 	a_8;
input 	a_9;
input 	a_10;
input 	a_11;
input 	a_12;
output 	dffe18;
output 	dffe17;
output 	dffe15;
output 	dffe16;
output 	dffe1;
output 	dffe2;
output 	dffe3;
output 	dffe4;
output 	dffe5;
output 	dffe6;
output 	dffe7;
output 	dffe8;
output 	dffe9;
output 	dffe10;
output 	dffe11;
output 	dffe12;
output 	dffe13;
output 	dffe14;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_add_sub_jdg_10 auto_generated(
	.a_17(a_17),
	.xordvalue_10(xordvalue_10),
	.a_16(a_16),
	.a_15(a_15),
	.a_14(a_14),
	.a_13(a_13),
	.a_0(a_0),
	.xordvalue_0(xordvalue_0),
	.a_1(a_1),
	.xordvalue_1(xordvalue_1),
	.a_2(a_2),
	.xordvalue_2(xordvalue_2),
	.a_3(a_3),
	.xordvalue_3(xordvalue_3),
	.a_4(a_4),
	.a_5(a_5),
	.a_6(a_6),
	.a_7(a_7),
	.a_8(a_8),
	.a_9(a_9),
	.a_10(a_10),
	.a_11(a_11),
	.a_12(a_12),
	.dffe181(dffe18),
	.dffe171(dffe17),
	.dffe151(dffe15),
	.dffe161(dffe16),
	.dffe19(dffe1),
	.dffe21(dffe2),
	.dffe31(dffe3),
	.dffe41(dffe4),
	.dffe51(dffe5),
	.dffe61(dffe6),
	.dffe71(dffe7),
	.dffe81(dffe8),
	.dffe91(dffe9),
	.dffe101(dffe10),
	.dffe111(dffe11),
	.dffe121(dffe12),
	.dffe131(dffe13),
	.dffe141(dffe14),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module nco_test_add_sub_jdg_10 (
	a_17,
	xordvalue_10,
	a_16,
	a_15,
	a_14,
	a_13,
	a_0,
	xordvalue_0,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	xordvalue_3,
	a_4,
	a_5,
	a_6,
	a_7,
	a_8,
	a_9,
	a_10,
	a_11,
	a_12,
	dffe181,
	dffe171,
	dffe151,
	dffe161,
	dffe19,
	dffe21,
	dffe31,
	dffe41,
	dffe51,
	dffe61,
	dffe71,
	dffe81,
	dffe91,
	dffe101,
	dffe111,
	dffe121,
	dffe131,
	dffe141,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_10;
input 	a_16;
input 	a_15;
input 	a_14;
input 	a_13;
input 	a_0;
input 	xordvalue_0;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	xordvalue_3;
input 	a_4;
input 	a_5;
input 	a_6;
input 	a_7;
input 	a_8;
input 	a_9;
input 	a_10;
input 	a_11;
input 	a_12;
output 	dffe181;
output 	dffe171;
output 	dffe151;
output 	dffe161;
output 	dffe19;
output 	dffe21;
output 	dffe31;
output 	dffe41;
output 	dffe51;
output 	dffe61;
output 	dffe71;
output 	dffe81;
output 	dffe91;
output 	dffe101;
output 	dffe111;
output 	dffe121;
output 	dffe131;
output 	dffe141;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~COUT ;
wire \add_sub_cella[12]~COUT ;
wire \add_sub_cella[13]~COUT ;
wire \add_sub_cella[14]~COUT ;
wire \add_sub_cella[15]~COUT ;
wire \add_sub_cella[16]~COUT ;
wire \add_sub_cella[17]~sumout ;
wire \add_sub_cella[16]~sumout ;
wire \add_sub_cella[14]~sumout ;
wire \add_sub_cella[15]~sumout ;
wire \add_sub_cella[0]~sumout ;
wire \add_sub_cella[1]~sumout ;
wire \add_sub_cella[2]~sumout ;
wire \add_sub_cella[3]~sumout ;
wire \add_sub_cella[4]~sumout ;
wire \add_sub_cella[5]~sumout ;
wire \add_sub_cella[6]~sumout ;
wire \add_sub_cella[7]~sumout ;
wire \add_sub_cella[8]~sumout ;
wire \add_sub_cella[9]~sumout ;
wire \add_sub_cella[10]~sumout ;
wire \add_sub_cella[11]~sumout ;
wire \add_sub_cella[12]~sumout ;
wire \add_sub_cella[13]~sumout ;


dffeas dffe18(
	.clk(clock),
	.d(\add_sub_cella[17]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe181),
	.prn(vcc));
defparam dffe18.is_wysiwyg = "true";
defparam dffe18.power_up = "low";

dffeas dffe17(
	.clk(clock),
	.d(\add_sub_cella[16]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe171),
	.prn(vcc));
defparam dffe17.is_wysiwyg = "true";
defparam dffe17.power_up = "low";

dffeas dffe15(
	.clk(clock),
	.d(\add_sub_cella[14]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe151),
	.prn(vcc));
defparam dffe15.is_wysiwyg = "true";
defparam dffe15.power_up = "low";

dffeas dffe16(
	.clk(clock),
	.d(\add_sub_cella[15]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe161),
	.prn(vcc));
defparam dffe16.is_wysiwyg = "true";
defparam dffe16.power_up = "low";

dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe19),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

dffeas dffe13(
	.clk(clock),
	.d(\add_sub_cella[12]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe131),
	.prn(vcc));
defparam dffe13.is_wysiwyg = "true";
defparam dffe13.power_up = "low";

dffeas dffe14(
	.clk(clock),
	.d(\add_sub_cella[13]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe141),
	.prn(vcc));
defparam dffe14.is_wysiwyg = "true";
defparam dffe14.power_up = "low";

arriav_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_1),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_2),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_3),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(\add_sub_cella[11]~COUT ),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[12] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[11]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[12]~sumout ),
	.cout(\add_sub_cella[12]~COUT ),
	.shareout());
defparam \add_sub_cella[12] .extended_lut = "off";
defparam \add_sub_cella[12] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[12] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[13] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[12]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[13]~sumout ),
	.cout(\add_sub_cella[13]~COUT ),
	.shareout());
defparam \add_sub_cella[13] .extended_lut = "off";
defparam \add_sub_cella[13] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[13] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[14] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[13]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[14]~sumout ),
	.cout(\add_sub_cella[14]~COUT ),
	.shareout());
defparam \add_sub_cella[14] .extended_lut = "off";
defparam \add_sub_cella[14] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[14] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[15] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[14]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[15]~sumout ),
	.cout(\add_sub_cella[15]~COUT ),
	.shareout());
defparam \add_sub_cella[15] .extended_lut = "off";
defparam \add_sub_cella[15] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[15] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[16] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_16),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[15]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[16]~sumout ),
	.cout(\add_sub_cella[16]~COUT ),
	.shareout());
defparam \add_sub_cella[16] .extended_lut = "off";
defparam \add_sub_cella[16] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[16] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[17] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_17),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[16]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[17]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[17] .extended_lut = "off";
defparam \add_sub_cella[17] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[17] .shared_arith = "off";

endmodule

module nco_test_cordic_sxor_1p_lpm_12 (
	sin_o_0,
	dffe18,
	dffe16,
	dffe17,
	dffe161,
	pipeline_dffe_17,
	dffe1,
	dffe181,
	dffe2,
	dffe3,
	dffe4,
	dffe5,
	dffe6,
	dffe7,
	dffe8,
	dffe9,
	dffe10,
	dffe11,
	dffe12,
	dffe13,
	dffe14,
	dffe15,
	dffe171,
	pipeline_dffe_16,
	dffe151,
	dffe162,
	pipeline_dffe_14,
	pipeline_dffe_15,
	dffe19,
	dffe21,
	dffe31,
	dffe41,
	dffe51,
	dffe61,
	dffe71,
	dffe81,
	dffe91,
	dffe101,
	dffe111,
	dffe121,
	dffe131,
	dffe141,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	sin_o_0;
output 	dffe18;
output 	dffe16;
output 	dffe17;
input 	dffe161;
input 	pipeline_dffe_17;
output 	dffe1;
input 	dffe181;
output 	dffe2;
output 	dffe3;
output 	dffe4;
output 	dffe5;
output 	dffe6;
output 	dffe7;
output 	dffe8;
output 	dffe9;
output 	dffe10;
output 	dffe11;
output 	dffe12;
output 	dffe13;
output 	dffe14;
output 	dffe15;
input 	dffe171;
input 	pipeline_dffe_16;
input 	dffe151;
input 	dffe162;
input 	pipeline_dffe_14;
input 	pipeline_dffe_15;
input 	dffe19;
input 	dffe21;
input 	dffe31;
input 	dffe41;
input 	dffe51;
input 	dffe61;
input 	dffe71;
input 	dffe81;
input 	dffe91;
input 	dffe101;
input 	dffe111;
input 	dffe121;
input 	dffe131;
input 	dffe141;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[17]~q ;
wire \xordvalue[10]~q ;
wire \Add0~1_sumout ;
wire \a[16]~q ;
wire \a[15]~q ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \a[14]~q ;
wire \a[0]~q ;
wire \xordvalue[0]~q ;
wire \a[1]~q ;
wire \xordvalue[1]~q ;
wire \a[2]~q ;
wire \xordvalue[2]~q ;
wire \a[3]~q ;
wire \a[4]~q ;
wire \a[5]~q ;
wire \a[6]~q ;
wire \a[7]~q ;
wire \a[8]~q ;
wire \a[9]~q ;
wire \a[10]~q ;
wire \a[11]~q ;
wire \a[12]~q ;
wire \a[13]~q ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~51 ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~55 ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~59 ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~63 ;
wire \Add0~65_sumout ;
wire \Add0~66 ;
wire \Add0~67 ;
wire \Add0~69_sumout ;
wire \Add0~70 ;
wire \Add0~71 ;
wire \xordvalue~0_combout ;
wire \xordvalue~1_combout ;
wire \xordvalue~2_combout ;
wire \xordvalue~3_combout ;


nco_test_lpm_add_sub_30 u0(
	.a_17(\a[17]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.a_16(\a[16]~q ),
	.a_15(\a[15]~q ),
	.a_14(\a[14]~q ),
	.a_0(\a[0]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_1(\a[1]~q ),
	.xordvalue_1(\xordvalue[1]~q ),
	.a_2(\a[2]~q ),
	.xordvalue_2(\xordvalue[2]~q ),
	.a_3(\a[3]~q ),
	.a_4(\a[4]~q ),
	.a_5(\a[5]~q ),
	.a_6(\a[6]~q ),
	.a_7(\a[7]~q ),
	.a_8(\a[8]~q ),
	.a_9(\a[9]~q ),
	.a_10(\a[10]~q ),
	.a_11(\a[11]~q ),
	.a_12(\a[12]~q ),
	.a_13(\a[13]~q ),
	.dffe18(dffe18),
	.dffe16(dffe16),
	.dffe17(dffe17),
	.dffe1(dffe1),
	.dffe2(dffe2),
	.dffe3(dffe3),
	.dffe4(dffe4),
	.dffe5(dffe5),
	.dffe6(dffe6),
	.dffe7(dffe7),
	.dffe8(dffe8),
	.dffe9(dffe9),
	.dffe10(dffe10),
	.dffe11(dffe11),
	.dffe12(dffe12),
	.dffe13(dffe13),
	.dffe14(dffe14),
	.dffe15(dffe15),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[17] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[17]~q ),
	.prn(vcc));
defparam \a[17] .is_wysiwyg = "true";
defparam \a[17] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe181),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "on";

dffeas \a[16] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[16]~q ),
	.prn(vcc));
defparam \a[16] .is_wysiwyg = "true";
defparam \a[16] .power_up = "low";

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe171),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~5 .shared_arith = "on";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe162),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~9 .shared_arith = "on";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \xordvalue[1] (
	.clk(clk),
	.d(\xordvalue~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[1]~q ),
	.prn(vcc));
defparam \xordvalue[1] .is_wysiwyg = "true";
defparam \xordvalue[1] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \xordvalue[2] (
	.clk(clk),
	.d(\xordvalue~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[2]~q ),
	.prn(vcc));
defparam \xordvalue[2] .is_wysiwyg = "true";
defparam \xordvalue[2] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~70 ),
	.sharein(\Add0~71 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~13 .shared_arith = "on";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!dffe19),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add0~17 .shared_arith = "on";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "on";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~25 .shared_arith = "on";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~29 .shared_arith = "on";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~33 .shared_arith = "on";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~37 .shared_arith = "on";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~41 .shared_arith = "on";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout(\Add0~47 ));
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~45 .shared_arith = "on";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(\Add0~47 ),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout(\Add0~51 ));
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~49 .shared_arith = "on";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(\Add0~51 ),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout(\Add0~55 ));
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~53 .shared_arith = "on";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(\Add0~55 ),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout(\Add0~59 ));
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~57 .shared_arith = "on";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(\Add0~59 ),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout(\Add0~63 ));
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~61 .shared_arith = "on";

arriav_lcell_comb \Add0~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(\Add0~63 ),
	.combout(),
	.sumout(\Add0~65_sumout ),
	.cout(\Add0~66 ),
	.shareout(\Add0~67 ));
defparam \Add0~65 .extended_lut = "off";
defparam \Add0~65 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~65 .shared_arith = "on";

arriav_lcell_comb \Add0~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~66 ),
	.sharein(\Add0~67 ),
	.combout(),
	.sumout(\Add0~69_sumout ),
	.cout(\Add0~70 ),
	.shareout(\Add0~71 ));
defparam \Add0~69 .extended_lut = "off";
defparam \Add0~69 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~69 .shared_arith = "on";

arriav_lcell_comb \xordvalue~0 (
	.dataa(!dffe161),
	.datab(!pipeline_dffe_17),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

arriav_lcell_comb \xordvalue~1 (
	.dataa(!dffe161),
	.datab(!pipeline_dffe_14),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~1 .extended_lut = "off";
defparam \xordvalue~1 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~1 .shared_arith = "off";

arriav_lcell_comb \xordvalue~2 (
	.dataa(!dffe161),
	.datab(!pipeline_dffe_15),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~2 .extended_lut = "off";
defparam \xordvalue~2 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~2 .shared_arith = "off";

arriav_lcell_comb \xordvalue~3 (
	.dataa(!dffe161),
	.datab(!pipeline_dffe_16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~3 .extended_lut = "off";
defparam \xordvalue~3 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~3 .shared_arith = "off";

endmodule

module nco_test_lpm_add_sub_30 (
	a_17,
	xordvalue_10,
	a_16,
	a_15,
	a_14,
	a_0,
	xordvalue_0,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	a_4,
	a_5,
	a_6,
	a_7,
	a_8,
	a_9,
	a_10,
	a_11,
	a_12,
	a_13,
	dffe18,
	dffe16,
	dffe17,
	dffe1,
	dffe2,
	dffe3,
	dffe4,
	dffe5,
	dffe6,
	dffe7,
	dffe8,
	dffe9,
	dffe10,
	dffe11,
	dffe12,
	dffe13,
	dffe14,
	dffe15,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_10;
input 	a_16;
input 	a_15;
input 	a_14;
input 	a_0;
input 	xordvalue_0;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	a_4;
input 	a_5;
input 	a_6;
input 	a_7;
input 	a_8;
input 	a_9;
input 	a_10;
input 	a_11;
input 	a_12;
input 	a_13;
output 	dffe18;
output 	dffe16;
output 	dffe17;
output 	dffe1;
output 	dffe2;
output 	dffe3;
output 	dffe4;
output 	dffe5;
output 	dffe6;
output 	dffe7;
output 	dffe8;
output 	dffe9;
output 	dffe10;
output 	dffe11;
output 	dffe12;
output 	dffe13;
output 	dffe14;
output 	dffe15;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_add_sub_jdg_11 auto_generated(
	.a_17(a_17),
	.xordvalue_10(xordvalue_10),
	.a_16(a_16),
	.a_15(a_15),
	.a_14(a_14),
	.a_0(a_0),
	.xordvalue_0(xordvalue_0),
	.a_1(a_1),
	.xordvalue_1(xordvalue_1),
	.a_2(a_2),
	.xordvalue_2(xordvalue_2),
	.a_3(a_3),
	.a_4(a_4),
	.a_5(a_5),
	.a_6(a_6),
	.a_7(a_7),
	.a_8(a_8),
	.a_9(a_9),
	.a_10(a_10),
	.a_11(a_11),
	.a_12(a_12),
	.a_13(a_13),
	.dffe181(dffe18),
	.dffe161(dffe16),
	.dffe171(dffe17),
	.dffe19(dffe1),
	.dffe21(dffe2),
	.dffe31(dffe3),
	.dffe41(dffe4),
	.dffe51(dffe5),
	.dffe61(dffe6),
	.dffe71(dffe7),
	.dffe81(dffe8),
	.dffe91(dffe9),
	.dffe101(dffe10),
	.dffe111(dffe11),
	.dffe121(dffe12),
	.dffe131(dffe13),
	.dffe141(dffe14),
	.dffe151(dffe15),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module nco_test_add_sub_jdg_11 (
	a_17,
	xordvalue_10,
	a_16,
	a_15,
	a_14,
	a_0,
	xordvalue_0,
	a_1,
	xordvalue_1,
	a_2,
	xordvalue_2,
	a_3,
	a_4,
	a_5,
	a_6,
	a_7,
	a_8,
	a_9,
	a_10,
	a_11,
	a_12,
	a_13,
	dffe181,
	dffe161,
	dffe171,
	dffe19,
	dffe21,
	dffe31,
	dffe41,
	dffe51,
	dffe61,
	dffe71,
	dffe81,
	dffe91,
	dffe101,
	dffe111,
	dffe121,
	dffe131,
	dffe141,
	dffe151,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_10;
input 	a_16;
input 	a_15;
input 	a_14;
input 	a_0;
input 	xordvalue_0;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	xordvalue_2;
input 	a_3;
input 	a_4;
input 	a_5;
input 	a_6;
input 	a_7;
input 	a_8;
input 	a_9;
input 	a_10;
input 	a_11;
input 	a_12;
input 	a_13;
output 	dffe181;
output 	dffe161;
output 	dffe171;
output 	dffe19;
output 	dffe21;
output 	dffe31;
output 	dffe41;
output 	dffe51;
output 	dffe61;
output 	dffe71;
output 	dffe81;
output 	dffe91;
output 	dffe101;
output 	dffe111;
output 	dffe121;
output 	dffe131;
output 	dffe141;
output 	dffe151;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~COUT ;
wire \add_sub_cella[12]~COUT ;
wire \add_sub_cella[13]~COUT ;
wire \add_sub_cella[14]~COUT ;
wire \add_sub_cella[15]~COUT ;
wire \add_sub_cella[16]~COUT ;
wire \add_sub_cella[17]~sumout ;
wire \add_sub_cella[15]~sumout ;
wire \add_sub_cella[16]~sumout ;
wire \add_sub_cella[0]~sumout ;
wire \add_sub_cella[1]~sumout ;
wire \add_sub_cella[2]~sumout ;
wire \add_sub_cella[3]~sumout ;
wire \add_sub_cella[4]~sumout ;
wire \add_sub_cella[5]~sumout ;
wire \add_sub_cella[6]~sumout ;
wire \add_sub_cella[7]~sumout ;
wire \add_sub_cella[8]~sumout ;
wire \add_sub_cella[9]~sumout ;
wire \add_sub_cella[10]~sumout ;
wire \add_sub_cella[11]~sumout ;
wire \add_sub_cella[12]~sumout ;
wire \add_sub_cella[13]~sumout ;
wire \add_sub_cella[14]~sumout ;


dffeas dffe18(
	.clk(clock),
	.d(\add_sub_cella[17]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe181),
	.prn(vcc));
defparam dffe18.is_wysiwyg = "true";
defparam dffe18.power_up = "low";

dffeas dffe16(
	.clk(clock),
	.d(\add_sub_cella[15]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe161),
	.prn(vcc));
defparam dffe16.is_wysiwyg = "true";
defparam dffe16.power_up = "low";

dffeas dffe17(
	.clk(clock),
	.d(\add_sub_cella[16]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe171),
	.prn(vcc));
defparam dffe17.is_wysiwyg = "true";
defparam dffe17.power_up = "low";

dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe19),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

dffeas dffe13(
	.clk(clock),
	.d(\add_sub_cella[12]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe131),
	.prn(vcc));
defparam dffe13.is_wysiwyg = "true";
defparam dffe13.power_up = "low";

dffeas dffe14(
	.clk(clock),
	.d(\add_sub_cella[13]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe141),
	.prn(vcc));
defparam dffe14.is_wysiwyg = "true";
defparam dffe14.power_up = "low";

dffeas dffe15(
	.clk(clock),
	.d(\add_sub_cella[14]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe151),
	.prn(vcc));
defparam dffe15.is_wysiwyg = "true";
defparam dffe15.power_up = "low";

arriav_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_1),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_2),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(\add_sub_cella[11]~COUT ),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[12] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[11]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[12]~sumout ),
	.cout(\add_sub_cella[12]~COUT ),
	.shareout());
defparam \add_sub_cella[12] .extended_lut = "off";
defparam \add_sub_cella[12] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[12] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[13] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[12]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[13]~sumout ),
	.cout(\add_sub_cella[13]~COUT ),
	.shareout());
defparam \add_sub_cella[13] .extended_lut = "off";
defparam \add_sub_cella[13] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[13] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[14] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[13]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[14]~sumout ),
	.cout(\add_sub_cella[14]~COUT ),
	.shareout());
defparam \add_sub_cella[14] .extended_lut = "off";
defparam \add_sub_cella[14] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[14] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[15] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[14]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[15]~sumout ),
	.cout(\add_sub_cella[15]~COUT ),
	.shareout());
defparam \add_sub_cella[15] .extended_lut = "off";
defparam \add_sub_cella[15] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[15] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[16] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_16),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[15]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[16]~sumout ),
	.cout(\add_sub_cella[16]~COUT ),
	.shareout());
defparam \add_sub_cella[16] .extended_lut = "off";
defparam \add_sub_cella[16] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[16] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[17] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_17),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[16]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[17]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[17] .extended_lut = "off";
defparam \add_sub_cella[17] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[17] .shared_arith = "off";

endmodule

module nco_test_cordic_sxor_1p_lpm_13 (
	sin_o_0,
	dffe18,
	dffe17,
	dffe1,
	dffe2,
	dffe3,
	dffe4,
	dffe5,
	dffe6,
	dffe7,
	dffe8,
	dffe9,
	dffe10,
	dffe11,
	dffe12,
	dffe13,
	dffe14,
	dffe15,
	dffe16,
	dffe161,
	dffe181,
	pipeline_dffe_17,
	dffe162,
	dffe171,
	pipeline_dffe_16,
	pipeline_dffe_15,
	dffe19,
	dffe21,
	dffe31,
	dffe41,
	dffe51,
	dffe61,
	dffe71,
	dffe81,
	dffe91,
	dffe101,
	dffe111,
	dffe121,
	dffe131,
	dffe141,
	dffe151,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	sin_o_0;
output 	dffe18;
output 	dffe17;
output 	dffe1;
output 	dffe2;
output 	dffe3;
output 	dffe4;
output 	dffe5;
output 	dffe6;
output 	dffe7;
output 	dffe8;
output 	dffe9;
output 	dffe10;
output 	dffe11;
output 	dffe12;
output 	dffe13;
output 	dffe14;
output 	dffe15;
output 	dffe16;
input 	dffe161;
input 	dffe181;
input 	pipeline_dffe_17;
input 	dffe162;
input 	dffe171;
input 	pipeline_dffe_16;
input 	pipeline_dffe_15;
input 	dffe19;
input 	dffe21;
input 	dffe31;
input 	dffe41;
input 	dffe51;
input 	dffe61;
input 	dffe71;
input 	dffe81;
input 	dffe91;
input 	dffe101;
input 	dffe111;
input 	dffe121;
input 	dffe131;
input 	dffe141;
input 	dffe151;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[17]~q ;
wire \xordvalue[10]~q ;
wire \a[16]~q ;
wire \Add0~1_sumout ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \a[15]~q ;
wire \a[0]~q ;
wire \xordvalue[0]~q ;
wire \a[1]~q ;
wire \xordvalue[1]~q ;
wire \a[2]~q ;
wire \a[3]~q ;
wire \a[4]~q ;
wire \a[5]~q ;
wire \a[6]~q ;
wire \a[7]~q ;
wire \a[8]~q ;
wire \a[9]~q ;
wire \a[10]~q ;
wire \a[11]~q ;
wire \a[12]~q ;
wire \a[13]~q ;
wire \a[14]~q ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~51 ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~55 ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~59 ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~63 ;
wire \Add0~65_sumout ;
wire \Add0~66 ;
wire \Add0~67 ;
wire \Add0~69_sumout ;
wire \Add0~70 ;
wire \Add0~71 ;
wire \xordvalue~0_combout ;
wire \xordvalue~1_combout ;
wire \xordvalue~2_combout ;


nco_test_lpm_add_sub_31 u0(
	.a_17(\a[17]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.a_16(\a[16]~q ),
	.a_15(\a[15]~q ),
	.a_0(\a[0]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_1(\a[1]~q ),
	.xordvalue_1(\xordvalue[1]~q ),
	.a_2(\a[2]~q ),
	.a_3(\a[3]~q ),
	.a_4(\a[4]~q ),
	.a_5(\a[5]~q ),
	.a_6(\a[6]~q ),
	.a_7(\a[7]~q ),
	.a_8(\a[8]~q ),
	.a_9(\a[9]~q ),
	.a_10(\a[10]~q ),
	.a_11(\a[11]~q ),
	.a_12(\a[12]~q ),
	.a_13(\a[13]~q ),
	.a_14(\a[14]~q ),
	.dffe18(dffe18),
	.dffe17(dffe17),
	.dffe1(dffe1),
	.dffe2(dffe2),
	.dffe3(dffe3),
	.dffe4(dffe4),
	.dffe5(dffe5),
	.dffe6(dffe6),
	.dffe7(dffe7),
	.dffe8(dffe8),
	.dffe9(dffe9),
	.dffe10(dffe10),
	.dffe11(dffe11),
	.dffe12(dffe12),
	.dffe13(dffe13),
	.dffe14(dffe14),
	.dffe15(dffe15),
	.dffe16(dffe16),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[17] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[17]~q ),
	.prn(vcc));
defparam \a[17] .is_wysiwyg = "true";
defparam \a[17] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

dffeas \a[16] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[16]~q ),
	.prn(vcc));
defparam \a[16] .is_wysiwyg = "true";
defparam \a[16] .power_up = "low";

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe181),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "on";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe171),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~5 .shared_arith = "on";

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \xordvalue[1] (
	.clk(clk),
	.d(\xordvalue~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[1]~q ),
	.prn(vcc));
defparam \xordvalue[1] .is_wysiwyg = "true";
defparam \xordvalue[1] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe162),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~70 ),
	.sharein(\Add0~71 ),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~9 .shared_arith = "on";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!dffe19),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add0~13 .shared_arith = "on";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~17 .shared_arith = "on";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "on";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~25 .shared_arith = "on";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~29 .shared_arith = "on";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~33 .shared_arith = "on";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~37 .shared_arith = "on";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~41 .shared_arith = "on";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout(\Add0~47 ));
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~45 .shared_arith = "on";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(\Add0~47 ),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout(\Add0~51 ));
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~49 .shared_arith = "on";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(\Add0~51 ),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout(\Add0~55 ));
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~53 .shared_arith = "on";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(\Add0~55 ),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout(\Add0~59 ));
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~57 .shared_arith = "on";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(\Add0~59 ),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout(\Add0~63 ));
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~61 .shared_arith = "on";

arriav_lcell_comb \Add0~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(\Add0~63 ),
	.combout(),
	.sumout(\Add0~65_sumout ),
	.cout(\Add0~66 ),
	.shareout(\Add0~67 ));
defparam \Add0~65 .extended_lut = "off";
defparam \Add0~65 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~65 .shared_arith = "on";

arriav_lcell_comb \Add0~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~66 ),
	.sharein(\Add0~67 ),
	.combout(),
	.sumout(\Add0~69_sumout ),
	.cout(\Add0~70 ),
	.shareout(\Add0~71 ));
defparam \Add0~69 .extended_lut = "off";
defparam \Add0~69 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~69 .shared_arith = "on";

arriav_lcell_comb \xordvalue~0 (
	.dataa(!pipeline_dffe_17),
	.datab(!dffe161),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

arriav_lcell_comb \xordvalue~1 (
	.dataa(!pipeline_dffe_15),
	.datab(!dffe161),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~1 .extended_lut = "off";
defparam \xordvalue~1 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~1 .shared_arith = "off";

arriav_lcell_comb \xordvalue~2 (
	.dataa(!pipeline_dffe_16),
	.datab(!dffe161),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~2 .extended_lut = "off";
defparam \xordvalue~2 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~2 .shared_arith = "off";

endmodule

module nco_test_lpm_add_sub_31 (
	a_17,
	xordvalue_10,
	a_16,
	a_15,
	a_0,
	xordvalue_0,
	a_1,
	xordvalue_1,
	a_2,
	a_3,
	a_4,
	a_5,
	a_6,
	a_7,
	a_8,
	a_9,
	a_10,
	a_11,
	a_12,
	a_13,
	a_14,
	dffe18,
	dffe17,
	dffe1,
	dffe2,
	dffe3,
	dffe4,
	dffe5,
	dffe6,
	dffe7,
	dffe8,
	dffe9,
	dffe10,
	dffe11,
	dffe12,
	dffe13,
	dffe14,
	dffe15,
	dffe16,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_10;
input 	a_16;
input 	a_15;
input 	a_0;
input 	xordvalue_0;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	a_3;
input 	a_4;
input 	a_5;
input 	a_6;
input 	a_7;
input 	a_8;
input 	a_9;
input 	a_10;
input 	a_11;
input 	a_12;
input 	a_13;
input 	a_14;
output 	dffe18;
output 	dffe17;
output 	dffe1;
output 	dffe2;
output 	dffe3;
output 	dffe4;
output 	dffe5;
output 	dffe6;
output 	dffe7;
output 	dffe8;
output 	dffe9;
output 	dffe10;
output 	dffe11;
output 	dffe12;
output 	dffe13;
output 	dffe14;
output 	dffe15;
output 	dffe16;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_add_sub_jdg_12 auto_generated(
	.a_17(a_17),
	.xordvalue_10(xordvalue_10),
	.a_16(a_16),
	.a_15(a_15),
	.a_0(a_0),
	.xordvalue_0(xordvalue_0),
	.a_1(a_1),
	.xordvalue_1(xordvalue_1),
	.a_2(a_2),
	.a_3(a_3),
	.a_4(a_4),
	.a_5(a_5),
	.a_6(a_6),
	.a_7(a_7),
	.a_8(a_8),
	.a_9(a_9),
	.a_10(a_10),
	.a_11(a_11),
	.a_12(a_12),
	.a_13(a_13),
	.a_14(a_14),
	.dffe181(dffe18),
	.dffe171(dffe17),
	.dffe19(dffe1),
	.dffe21(dffe2),
	.dffe31(dffe3),
	.dffe41(dffe4),
	.dffe51(dffe5),
	.dffe61(dffe6),
	.dffe71(dffe7),
	.dffe81(dffe8),
	.dffe91(dffe9),
	.dffe101(dffe10),
	.dffe111(dffe11),
	.dffe121(dffe12),
	.dffe131(dffe13),
	.dffe141(dffe14),
	.dffe151(dffe15),
	.dffe161(dffe16),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module nco_test_add_sub_jdg_12 (
	a_17,
	xordvalue_10,
	a_16,
	a_15,
	a_0,
	xordvalue_0,
	a_1,
	xordvalue_1,
	a_2,
	a_3,
	a_4,
	a_5,
	a_6,
	a_7,
	a_8,
	a_9,
	a_10,
	a_11,
	a_12,
	a_13,
	a_14,
	dffe181,
	dffe171,
	dffe19,
	dffe21,
	dffe31,
	dffe41,
	dffe51,
	dffe61,
	dffe71,
	dffe81,
	dffe91,
	dffe101,
	dffe111,
	dffe121,
	dffe131,
	dffe141,
	dffe151,
	dffe161,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_10;
input 	a_16;
input 	a_15;
input 	a_0;
input 	xordvalue_0;
input 	a_1;
input 	xordvalue_1;
input 	a_2;
input 	a_3;
input 	a_4;
input 	a_5;
input 	a_6;
input 	a_7;
input 	a_8;
input 	a_9;
input 	a_10;
input 	a_11;
input 	a_12;
input 	a_13;
input 	a_14;
output 	dffe181;
output 	dffe171;
output 	dffe19;
output 	dffe21;
output 	dffe31;
output 	dffe41;
output 	dffe51;
output 	dffe61;
output 	dffe71;
output 	dffe81;
output 	dffe91;
output 	dffe101;
output 	dffe111;
output 	dffe121;
output 	dffe131;
output 	dffe141;
output 	dffe151;
output 	dffe161;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~COUT ;
wire \add_sub_cella[12]~COUT ;
wire \add_sub_cella[13]~COUT ;
wire \add_sub_cella[14]~COUT ;
wire \add_sub_cella[15]~COUT ;
wire \add_sub_cella[16]~COUT ;
wire \add_sub_cella[17]~sumout ;
wire \add_sub_cella[16]~sumout ;
wire \add_sub_cella[0]~sumout ;
wire \add_sub_cella[1]~sumout ;
wire \add_sub_cella[2]~sumout ;
wire \add_sub_cella[3]~sumout ;
wire \add_sub_cella[4]~sumout ;
wire \add_sub_cella[5]~sumout ;
wire \add_sub_cella[6]~sumout ;
wire \add_sub_cella[7]~sumout ;
wire \add_sub_cella[8]~sumout ;
wire \add_sub_cella[9]~sumout ;
wire \add_sub_cella[10]~sumout ;
wire \add_sub_cella[11]~sumout ;
wire \add_sub_cella[12]~sumout ;
wire \add_sub_cella[13]~sumout ;
wire \add_sub_cella[14]~sumout ;
wire \add_sub_cella[15]~sumout ;


dffeas dffe18(
	.clk(clock),
	.d(\add_sub_cella[17]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe181),
	.prn(vcc));
defparam dffe18.is_wysiwyg = "true";
defparam dffe18.power_up = "low";

dffeas dffe17(
	.clk(clock),
	.d(\add_sub_cella[16]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe171),
	.prn(vcc));
defparam dffe17.is_wysiwyg = "true";
defparam dffe17.power_up = "low";

dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe19),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

dffeas dffe13(
	.clk(clock),
	.d(\add_sub_cella[12]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe131),
	.prn(vcc));
defparam dffe13.is_wysiwyg = "true";
defparam dffe13.power_up = "low";

dffeas dffe14(
	.clk(clock),
	.d(\add_sub_cella[13]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe141),
	.prn(vcc));
defparam dffe14.is_wysiwyg = "true";
defparam dffe14.power_up = "low";

dffeas dffe15(
	.clk(clock),
	.d(\add_sub_cella[14]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe151),
	.prn(vcc));
defparam dffe15.is_wysiwyg = "true";
defparam dffe15.power_up = "low";

dffeas dffe16(
	.clk(clock),
	.d(\add_sub_cella[15]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe161),
	.prn(vcc));
defparam dffe16.is_wysiwyg = "true";
defparam dffe16.power_up = "low";

arriav_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_1),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(\add_sub_cella[11]~COUT ),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[12] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[11]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[12]~sumout ),
	.cout(\add_sub_cella[12]~COUT ),
	.shareout());
defparam \add_sub_cella[12] .extended_lut = "off";
defparam \add_sub_cella[12] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[12] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[13] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[12]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[13]~sumout ),
	.cout(\add_sub_cella[13]~COUT ),
	.shareout());
defparam \add_sub_cella[13] .extended_lut = "off";
defparam \add_sub_cella[13] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[13] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[14] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[13]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[14]~sumout ),
	.cout(\add_sub_cella[14]~COUT ),
	.shareout());
defparam \add_sub_cella[14] .extended_lut = "off";
defparam \add_sub_cella[14] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[14] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[15] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[14]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[15]~sumout ),
	.cout(\add_sub_cella[15]~COUT ),
	.shareout());
defparam \add_sub_cella[15] .extended_lut = "off";
defparam \add_sub_cella[15] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[15] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[16] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_16),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[15]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[16]~sumout ),
	.cout(\add_sub_cella[16]~COUT ),
	.shareout());
defparam \add_sub_cella[16] .extended_lut = "off";
defparam \add_sub_cella[16] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[16] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[17] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_17),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[16]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[17]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[17] .extended_lut = "off";
defparam \add_sub_cella[17] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[17] .shared_arith = "off";

endmodule

module nco_test_cordic_sxor_1p_lpm_14 (
	sin_o_0,
	dffe18,
	dffe1,
	dffe2,
	dffe3,
	dffe4,
	dffe5,
	dffe6,
	dffe7,
	dffe8,
	dffe9,
	dffe10,
	dffe11,
	dffe12,
	dffe13,
	dffe14,
	dffe15,
	dffe16,
	dffe17,
	dffe161,
	pipeline_dffe_17,
	dffe181,
	dffe171,
	pipeline_dffe_16,
	dffe19,
	dffe21,
	dffe31,
	dffe41,
	dffe51,
	dffe61,
	dffe71,
	dffe81,
	dffe91,
	dffe101,
	dffe111,
	dffe121,
	dffe131,
	dffe141,
	dffe151,
	dffe162,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	sin_o_0;
output 	dffe18;
output 	dffe1;
output 	dffe2;
output 	dffe3;
output 	dffe4;
output 	dffe5;
output 	dffe6;
output 	dffe7;
output 	dffe8;
output 	dffe9;
output 	dffe10;
output 	dffe11;
output 	dffe12;
output 	dffe13;
output 	dffe14;
output 	dffe15;
output 	dffe16;
output 	dffe17;
input 	dffe161;
input 	pipeline_dffe_17;
input 	dffe181;
input 	dffe171;
input 	pipeline_dffe_16;
input 	dffe19;
input 	dffe21;
input 	dffe31;
input 	dffe41;
input 	dffe51;
input 	dffe61;
input 	dffe71;
input 	dffe81;
input 	dffe91;
input 	dffe101;
input 	dffe111;
input 	dffe121;
input 	dffe131;
input 	dffe141;
input 	dffe151;
input 	dffe162;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[17]~q ;
wire \xordvalue[10]~q ;
wire \Add0~1_sumout ;
wire \a[16]~q ;
wire \a[0]~q ;
wire \xordvalue[0]~q ;
wire \a[1]~q ;
wire \a[2]~q ;
wire \a[3]~q ;
wire \a[4]~q ;
wire \a[5]~q ;
wire \a[6]~q ;
wire \a[7]~q ;
wire \a[8]~q ;
wire \a[9]~q ;
wire \a[10]~q ;
wire \a[11]~q ;
wire \a[12]~q ;
wire \a[13]~q ;
wire \a[14]~q ;
wire \a[15]~q ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~51 ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~55 ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~59 ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~63 ;
wire \Add0~65_sumout ;
wire \Add0~66 ;
wire \Add0~67 ;
wire \Add0~69_sumout ;
wire \Add0~70 ;
wire \Add0~71 ;
wire \xordvalue~0_combout ;
wire \xordvalue~1_combout ;


nco_test_lpm_add_sub_32 u0(
	.a_17(\a[17]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.a_16(\a[16]~q ),
	.a_0(\a[0]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_1(\a[1]~q ),
	.a_2(\a[2]~q ),
	.a_3(\a[3]~q ),
	.a_4(\a[4]~q ),
	.a_5(\a[5]~q ),
	.a_6(\a[6]~q ),
	.a_7(\a[7]~q ),
	.a_8(\a[8]~q ),
	.a_9(\a[9]~q ),
	.a_10(\a[10]~q ),
	.a_11(\a[11]~q ),
	.a_12(\a[12]~q ),
	.a_13(\a[13]~q ),
	.a_14(\a[14]~q ),
	.a_15(\a[15]~q ),
	.dffe18(dffe18),
	.dffe1(dffe1),
	.dffe2(dffe2),
	.dffe3(dffe3),
	.dffe4(dffe4),
	.dffe5(dffe5),
	.dffe6(dffe6),
	.dffe7(dffe7),
	.dffe8(dffe8),
	.dffe9(dffe9),
	.dffe10(dffe10),
	.dffe11(dffe11),
	.dffe12(dffe12),
	.dffe13(dffe13),
	.dffe14(dffe14),
	.dffe15(dffe15),
	.dffe16(dffe16),
	.dffe17(dffe17),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[17] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[17]~q ),
	.prn(vcc));
defparam \a[17] .is_wysiwyg = "true";
defparam \a[17] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe181),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "on";

dffeas \a[16] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[16]~q ),
	.prn(vcc));
defparam \a[16] .is_wysiwyg = "true";
defparam \a[16] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe171),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~70 ),
	.sharein(\Add0~71 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~5 .shared_arith = "on";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!dffe19),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add0~9 .shared_arith = "on";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~13 .shared_arith = "on";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~17 .shared_arith = "on";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "on";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~25 .shared_arith = "on";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~29 .shared_arith = "on";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~33 .shared_arith = "on";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~37 .shared_arith = "on";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~41 .shared_arith = "on";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout(\Add0~47 ));
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~45 .shared_arith = "on";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(\Add0~47 ),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout(\Add0~51 ));
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~49 .shared_arith = "on";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(\Add0~51 ),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout(\Add0~55 ));
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~53 .shared_arith = "on";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(\Add0~55 ),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout(\Add0~59 ));
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~57 .shared_arith = "on";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(\Add0~59 ),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout(\Add0~63 ));
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~61 .shared_arith = "on";

arriav_lcell_comb \Add0~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(\Add0~63 ),
	.combout(),
	.sumout(\Add0~65_sumout ),
	.cout(\Add0~66 ),
	.shareout(\Add0~67 ));
defparam \Add0~65 .extended_lut = "off";
defparam \Add0~65 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~65 .shared_arith = "on";

arriav_lcell_comb \Add0~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe162),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~66 ),
	.sharein(\Add0~67 ),
	.combout(),
	.sumout(\Add0~69_sumout ),
	.cout(\Add0~70 ),
	.shareout(\Add0~71 ));
defparam \Add0~69 .extended_lut = "off";
defparam \Add0~69 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~69 .shared_arith = "on";

arriav_lcell_comb \xordvalue~0 (
	.dataa(!dffe161),
	.datab(!pipeline_dffe_17),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

arriav_lcell_comb \xordvalue~1 (
	.dataa(!dffe161),
	.datab(!pipeline_dffe_16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~1 .extended_lut = "off";
defparam \xordvalue~1 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~1 .shared_arith = "off";

endmodule

module nco_test_lpm_add_sub_32 (
	a_17,
	xordvalue_10,
	a_16,
	a_0,
	xordvalue_0,
	a_1,
	a_2,
	a_3,
	a_4,
	a_5,
	a_6,
	a_7,
	a_8,
	a_9,
	a_10,
	a_11,
	a_12,
	a_13,
	a_14,
	a_15,
	dffe18,
	dffe1,
	dffe2,
	dffe3,
	dffe4,
	dffe5,
	dffe6,
	dffe7,
	dffe8,
	dffe9,
	dffe10,
	dffe11,
	dffe12,
	dffe13,
	dffe14,
	dffe15,
	dffe16,
	dffe17,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_10;
input 	a_16;
input 	a_0;
input 	xordvalue_0;
input 	a_1;
input 	a_2;
input 	a_3;
input 	a_4;
input 	a_5;
input 	a_6;
input 	a_7;
input 	a_8;
input 	a_9;
input 	a_10;
input 	a_11;
input 	a_12;
input 	a_13;
input 	a_14;
input 	a_15;
output 	dffe18;
output 	dffe1;
output 	dffe2;
output 	dffe3;
output 	dffe4;
output 	dffe5;
output 	dffe6;
output 	dffe7;
output 	dffe8;
output 	dffe9;
output 	dffe10;
output 	dffe11;
output 	dffe12;
output 	dffe13;
output 	dffe14;
output 	dffe15;
output 	dffe16;
output 	dffe17;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_add_sub_jdg_13 auto_generated(
	.a_17(a_17),
	.xordvalue_10(xordvalue_10),
	.a_16(a_16),
	.a_0(a_0),
	.xordvalue_0(xordvalue_0),
	.a_1(a_1),
	.a_2(a_2),
	.a_3(a_3),
	.a_4(a_4),
	.a_5(a_5),
	.a_6(a_6),
	.a_7(a_7),
	.a_8(a_8),
	.a_9(a_9),
	.a_10(a_10),
	.a_11(a_11),
	.a_12(a_12),
	.a_13(a_13),
	.a_14(a_14),
	.a_15(a_15),
	.dffe181(dffe18),
	.dffe19(dffe1),
	.dffe21(dffe2),
	.dffe31(dffe3),
	.dffe41(dffe4),
	.dffe51(dffe5),
	.dffe61(dffe6),
	.dffe71(dffe7),
	.dffe81(dffe8),
	.dffe91(dffe9),
	.dffe101(dffe10),
	.dffe111(dffe11),
	.dffe121(dffe12),
	.dffe131(dffe13),
	.dffe141(dffe14),
	.dffe151(dffe15),
	.dffe161(dffe16),
	.dffe171(dffe17),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module nco_test_add_sub_jdg_13 (
	a_17,
	xordvalue_10,
	a_16,
	a_0,
	xordvalue_0,
	a_1,
	a_2,
	a_3,
	a_4,
	a_5,
	a_6,
	a_7,
	a_8,
	a_9,
	a_10,
	a_11,
	a_12,
	a_13,
	a_14,
	a_15,
	dffe181,
	dffe19,
	dffe21,
	dffe31,
	dffe41,
	dffe51,
	dffe61,
	dffe71,
	dffe81,
	dffe91,
	dffe101,
	dffe111,
	dffe121,
	dffe131,
	dffe141,
	dffe151,
	dffe161,
	dffe171,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_10;
input 	a_16;
input 	a_0;
input 	xordvalue_0;
input 	a_1;
input 	a_2;
input 	a_3;
input 	a_4;
input 	a_5;
input 	a_6;
input 	a_7;
input 	a_8;
input 	a_9;
input 	a_10;
input 	a_11;
input 	a_12;
input 	a_13;
input 	a_14;
input 	a_15;
output 	dffe181;
output 	dffe19;
output 	dffe21;
output 	dffe31;
output 	dffe41;
output 	dffe51;
output 	dffe61;
output 	dffe71;
output 	dffe81;
output 	dffe91;
output 	dffe101;
output 	dffe111;
output 	dffe121;
output 	dffe131;
output 	dffe141;
output 	dffe151;
output 	dffe161;
output 	dffe171;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~COUT ;
wire \add_sub_cella[12]~COUT ;
wire \add_sub_cella[13]~COUT ;
wire \add_sub_cella[14]~COUT ;
wire \add_sub_cella[15]~COUT ;
wire \add_sub_cella[16]~COUT ;
wire \add_sub_cella[17]~sumout ;
wire \add_sub_cella[0]~sumout ;
wire \add_sub_cella[1]~sumout ;
wire \add_sub_cella[2]~sumout ;
wire \add_sub_cella[3]~sumout ;
wire \add_sub_cella[4]~sumout ;
wire \add_sub_cella[5]~sumout ;
wire \add_sub_cella[6]~sumout ;
wire \add_sub_cella[7]~sumout ;
wire \add_sub_cella[8]~sumout ;
wire \add_sub_cella[9]~sumout ;
wire \add_sub_cella[10]~sumout ;
wire \add_sub_cella[11]~sumout ;
wire \add_sub_cella[12]~sumout ;
wire \add_sub_cella[13]~sumout ;
wire \add_sub_cella[14]~sumout ;
wire \add_sub_cella[15]~sumout ;
wire \add_sub_cella[16]~sumout ;


dffeas dffe18(
	.clk(clock),
	.d(\add_sub_cella[17]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe181),
	.prn(vcc));
defparam dffe18.is_wysiwyg = "true";
defparam dffe18.power_up = "low";

dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe19),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

dffeas dffe13(
	.clk(clock),
	.d(\add_sub_cella[12]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe131),
	.prn(vcc));
defparam dffe13.is_wysiwyg = "true";
defparam dffe13.power_up = "low";

dffeas dffe14(
	.clk(clock),
	.d(\add_sub_cella[13]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe141),
	.prn(vcc));
defparam dffe14.is_wysiwyg = "true";
defparam dffe14.power_up = "low";

dffeas dffe15(
	.clk(clock),
	.d(\add_sub_cella[14]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe151),
	.prn(vcc));
defparam dffe15.is_wysiwyg = "true";
defparam dffe15.power_up = "low";

dffeas dffe16(
	.clk(clock),
	.d(\add_sub_cella[15]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe161),
	.prn(vcc));
defparam dffe16.is_wysiwyg = "true";
defparam dffe16.power_up = "low";

dffeas dffe17(
	.clk(clock),
	.d(\add_sub_cella[16]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe171),
	.prn(vcc));
defparam dffe17.is_wysiwyg = "true";
defparam dffe17.power_up = "low";

arriav_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(\add_sub_cella[11]~COUT ),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[12] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[11]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[12]~sumout ),
	.cout(\add_sub_cella[12]~COUT ),
	.shareout());
defparam \add_sub_cella[12] .extended_lut = "off";
defparam \add_sub_cella[12] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[12] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[13] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[12]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[13]~sumout ),
	.cout(\add_sub_cella[13]~COUT ),
	.shareout());
defparam \add_sub_cella[13] .extended_lut = "off";
defparam \add_sub_cella[13] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[13] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[14] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[13]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[14]~sumout ),
	.cout(\add_sub_cella[14]~COUT ),
	.shareout());
defparam \add_sub_cella[14] .extended_lut = "off";
defparam \add_sub_cella[14] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[14] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[15] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[14]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[15]~sumout ),
	.cout(\add_sub_cella[15]~COUT ),
	.shareout());
defparam \add_sub_cella[15] .extended_lut = "off";
defparam \add_sub_cella[15] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[15] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[16] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_16),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[15]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[16]~sumout ),
	.cout(\add_sub_cella[16]~COUT ),
	.shareout());
defparam \add_sub_cella[16] .extended_lut = "off";
defparam \add_sub_cella[16] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[16] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[17] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_17),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[16]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[17]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[17] .extended_lut = "off";
defparam \add_sub_cella[17] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[17] .shared_arith = "off";

endmodule

module nco_test_lpm_add_sub_33 (
	a_0,
	xordvalue_11,
	a_17,
	a_16,
	a_15,
	a_14,
	a_13,
	a_12,
	a_11,
	a_10,
	a_9,
	a_8,
	a_7,
	a_6,
	a_5,
	a_4,
	a_3,
	a_2,
	a_1,
	a_01,
	dffe18,
	dffe17,
	dffe16,
	dffe15,
	dffe14,
	dffe13,
	dffe12,
	dffe11,
	dffe10,
	dffe9,
	dffe8,
	dffe7,
	dffe6,
	dffe5,
	dffe3,
	dffe4,
	dffe1,
	dffe2,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_0;
input 	xordvalue_11;
input 	a_17;
input 	a_16;
input 	a_15;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_10;
input 	a_9;
input 	a_8;
input 	a_7;
input 	a_6;
input 	a_5;
input 	a_4;
input 	a_3;
input 	a_2;
input 	a_1;
input 	a_01;
output 	dffe18;
output 	dffe17;
output 	dffe16;
output 	dffe15;
output 	dffe14;
output 	dffe13;
output 	dffe12;
output 	dffe11;
output 	dffe10;
output 	dffe9;
output 	dffe8;
output 	dffe7;
output 	dffe6;
output 	dffe5;
output 	dffe3;
output 	dffe4;
output 	dffe1;
output 	dffe2;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_add_sub_jdg_14 auto_generated(
	.a_0(a_0),
	.xordvalue_11(xordvalue_11),
	.a_17(a_17),
	.a_16(a_16),
	.a_15(a_15),
	.a_14(a_14),
	.a_13(a_13),
	.a_12(a_12),
	.a_11(a_11),
	.a_10(a_10),
	.a_9(a_9),
	.a_8(a_8),
	.a_7(a_7),
	.a_6(a_6),
	.a_5(a_5),
	.a_4(a_4),
	.a_3(a_3),
	.a_2(a_2),
	.a_1(a_1),
	.a_01(a_01),
	.dffe181(dffe18),
	.dffe171(dffe17),
	.dffe161(dffe16),
	.dffe151(dffe15),
	.dffe141(dffe14),
	.dffe131(dffe13),
	.dffe121(dffe12),
	.dffe111(dffe11),
	.dffe101(dffe10),
	.dffe91(dffe9),
	.dffe81(dffe8),
	.dffe71(dffe7),
	.dffe61(dffe6),
	.dffe51(dffe5),
	.dffe31(dffe3),
	.dffe41(dffe4),
	.dffe19(dffe1),
	.dffe21(dffe2),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module nco_test_add_sub_jdg_14 (
	a_0,
	xordvalue_11,
	a_17,
	a_16,
	a_15,
	a_14,
	a_13,
	a_12,
	a_11,
	a_10,
	a_9,
	a_8,
	a_7,
	a_6,
	a_5,
	a_4,
	a_3,
	a_2,
	a_1,
	a_01,
	dffe181,
	dffe171,
	dffe161,
	dffe151,
	dffe141,
	dffe131,
	dffe121,
	dffe111,
	dffe101,
	dffe91,
	dffe81,
	dffe71,
	dffe61,
	dffe51,
	dffe31,
	dffe41,
	dffe19,
	dffe21,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_0;
input 	xordvalue_11;
input 	a_17;
input 	a_16;
input 	a_15;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_10;
input 	a_9;
input 	a_8;
input 	a_7;
input 	a_6;
input 	a_5;
input 	a_4;
input 	a_3;
input 	a_2;
input 	a_1;
input 	a_01;
output 	dffe181;
output 	dffe171;
output 	dffe161;
output 	dffe151;
output 	dffe141;
output 	dffe131;
output 	dffe121;
output 	dffe111;
output 	dffe101;
output 	dffe91;
output 	dffe81;
output 	dffe71;
output 	dffe61;
output 	dffe51;
output 	dffe31;
output 	dffe41;
output 	dffe19;
output 	dffe21;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~COUT ;
wire \add_sub_cella[12]~COUT ;
wire \add_sub_cella[13]~COUT ;
wire \add_sub_cella[14]~COUT ;
wire \add_sub_cella[15]~COUT ;
wire \add_sub_cella[16]~COUT ;
wire \add_sub_cella[17]~sumout ;
wire \add_sub_cella[16]~sumout ;
wire \add_sub_cella[15]~sumout ;
wire \add_sub_cella[14]~sumout ;
wire \add_sub_cella[13]~sumout ;
wire \add_sub_cella[12]~sumout ;
wire \add_sub_cella[11]~sumout ;
wire \add_sub_cella[10]~sumout ;
wire \add_sub_cella[9]~sumout ;
wire \add_sub_cella[8]~sumout ;
wire \add_sub_cella[7]~sumout ;
wire \add_sub_cella[6]~sumout ;
wire \add_sub_cella[5]~sumout ;
wire \add_sub_cella[4]~sumout ;
wire \add_sub_cella[2]~sumout ;
wire \add_sub_cella[3]~sumout ;
wire \add_sub_cella[0]~sumout ;
wire \add_sub_cella[1]~sumout ;


dffeas dffe18(
	.clk(clock),
	.d(\add_sub_cella[17]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe181),
	.prn(vcc));
defparam dffe18.is_wysiwyg = "true";
defparam dffe18.power_up = "low";

dffeas dffe17(
	.clk(clock),
	.d(\add_sub_cella[16]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe171),
	.prn(vcc));
defparam dffe17.is_wysiwyg = "true";
defparam dffe17.power_up = "low";

dffeas dffe16(
	.clk(clock),
	.d(\add_sub_cella[15]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe161),
	.prn(vcc));
defparam dffe16.is_wysiwyg = "true";
defparam dffe16.power_up = "low";

dffeas dffe15(
	.clk(clock),
	.d(\add_sub_cella[14]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe151),
	.prn(vcc));
defparam dffe15.is_wysiwyg = "true";
defparam dffe15.power_up = "low";

dffeas dffe14(
	.clk(clock),
	.d(\add_sub_cella[13]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe141),
	.prn(vcc));
defparam dffe14.is_wysiwyg = "true";
defparam dffe14.power_up = "low";

dffeas dffe13(
	.clk(clock),
	.d(\add_sub_cella[12]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe131),
	.prn(vcc));
defparam dffe13.is_wysiwyg = "true";
defparam dffe13.power_up = "low";

dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe19),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

arriav_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_01),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_11),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_11),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_11),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_11),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_11),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_11),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_11),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(\add_sub_cella[11]~COUT ),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[12] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_11),
	.datag(gnd),
	.cin(\add_sub_cella[11]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[12]~sumout ),
	.cout(\add_sub_cella[12]~COUT ),
	.shareout());
defparam \add_sub_cella[12] .extended_lut = "off";
defparam \add_sub_cella[12] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[12] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[13] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(\add_sub_cella[12]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[13]~sumout ),
	.cout(\add_sub_cella[13]~COUT ),
	.shareout());
defparam \add_sub_cella[13] .extended_lut = "off";
defparam \add_sub_cella[13] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[13] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[14] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(\add_sub_cella[13]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[14]~sumout ),
	.cout(\add_sub_cella[14]~COUT ),
	.shareout());
defparam \add_sub_cella[14] .extended_lut = "off";
defparam \add_sub_cella[14] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[14] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[15] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_11),
	.datag(gnd),
	.cin(\add_sub_cella[14]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[15]~sumout ),
	.cout(\add_sub_cella[15]~COUT ),
	.shareout());
defparam \add_sub_cella[15] .extended_lut = "off";
defparam \add_sub_cella[15] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[15] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[16] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_16),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(\add_sub_cella[15]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[16]~sumout ),
	.cout(\add_sub_cella[16]~COUT ),
	.shareout());
defparam \add_sub_cella[16] .extended_lut = "off";
defparam \add_sub_cella[16] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[16] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[17] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_17),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(\add_sub_cella[16]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[17]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[17] .extended_lut = "off";
defparam \add_sub_cella[17] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[17] .shared_arith = "off";

endmodule

module nco_test_cordic_sxor_1p_lpm_15 (
	sin_o_0,
	dffe1,
	dffe2,
	dffe3,
	dffe4,
	dffe5,
	dffe6,
	dffe7,
	dffe8,
	dffe9,
	dffe10,
	dffe11,
	dffe12,
	dffe13,
	dffe14,
	dffe15,
	dffe16,
	dffe17,
	dffe18,
	dffe161,
	dffe181,
	pipeline_dffe_17,
	dffe19,
	dffe21,
	dffe31,
	dffe41,
	dffe51,
	dffe61,
	dffe71,
	dffe81,
	dffe91,
	dffe101,
	dffe111,
	dffe121,
	dffe131,
	dffe141,
	dffe151,
	dffe162,
	dffe171,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	sin_o_0;
output 	dffe1;
output 	dffe2;
output 	dffe3;
output 	dffe4;
output 	dffe5;
output 	dffe6;
output 	dffe7;
output 	dffe8;
output 	dffe9;
output 	dffe10;
output 	dffe11;
output 	dffe12;
output 	dffe13;
output 	dffe14;
output 	dffe15;
output 	dffe16;
output 	dffe17;
output 	dffe18;
input 	dffe161;
input 	dffe181;
input 	pipeline_dffe_17;
input 	dffe19;
input 	dffe21;
input 	dffe31;
input 	dffe41;
input 	dffe51;
input 	dffe61;
input 	dffe71;
input 	dffe81;
input 	dffe91;
input 	dffe101;
input 	dffe111;
input 	dffe121;
input 	dffe131;
input 	dffe141;
input 	dffe151;
input 	dffe162;
input 	dffe171;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[0]~q ;
wire \xordvalue[0]~q ;
wire \a[1]~q ;
wire \a[2]~q ;
wire \a[3]~q ;
wire \a[4]~q ;
wire \a[5]~q ;
wire \a[6]~q ;
wire \a[7]~q ;
wire \a[8]~q ;
wire \a[9]~q ;
wire \a[10]~q ;
wire \a[11]~q ;
wire \a[12]~q ;
wire \a[13]~q ;
wire \a[14]~q ;
wire \a[15]~q ;
wire \a[16]~q ;
wire \a[17]~q ;
wire \Add0~1_sumout ;
wire \Add0~2 ;
wire \Add0~3 ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~51 ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~55 ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~59 ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~63 ;
wire \Add0~65_sumout ;
wire \Add0~66 ;
wire \Add0~67 ;
wire \Add0~69_sumout ;
wire \xordvalue~0_combout ;


nco_test_lpm_add_sub_34 u0(
	.a_0(\a[0]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_1(\a[1]~q ),
	.a_2(\a[2]~q ),
	.a_3(\a[3]~q ),
	.a_4(\a[4]~q ),
	.a_5(\a[5]~q ),
	.a_6(\a[6]~q ),
	.a_7(\a[7]~q ),
	.a_8(\a[8]~q ),
	.a_9(\a[9]~q ),
	.a_10(\a[10]~q ),
	.a_11(\a[11]~q ),
	.a_12(\a[12]~q ),
	.a_13(\a[13]~q ),
	.a_14(\a[14]~q ),
	.a_15(\a[15]~q ),
	.a_16(\a[16]~q ),
	.a_17(\a[17]~q ),
	.dffe1(dffe1),
	.dffe2(dffe2),
	.dffe3(dffe3),
	.dffe4(dffe4),
	.dffe5(dffe5),
	.dffe6(dffe6),
	.dffe7(dffe7),
	.dffe8(dffe8),
	.dffe9(dffe9),
	.dffe10(dffe10),
	.dffe11(dffe11),
	.dffe12(dffe12),
	.dffe13(dffe13),
	.dffe14(dffe14),
	.dffe15(dffe15),
	.dffe16(dffe16),
	.dffe17(dffe17),
	.dffe18(dffe18),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

dffeas \a[16] (
	.clk(clk),
	.d(\Add0~65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[16]~q ),
	.prn(vcc));
defparam \a[16] .is_wysiwyg = "true";
defparam \a[16] .power_up = "low";

dffeas \a[17] (
	.clk(clk),
	.d(\Add0~69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[17]~q ),
	.prn(vcc));
defparam \a[17] .is_wysiwyg = "true";
defparam \a[17] .power_up = "low";

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!dffe19),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(\Add0~2 ),
	.shareout(\Add0~3 ));
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add0~1 .shared_arith = "on";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~2 ),
	.sharein(\Add0~3 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~5 .shared_arith = "on";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~9 .shared_arith = "on";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~13 .shared_arith = "on";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~17 .shared_arith = "on";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "on";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~25 .shared_arith = "on";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~29 .shared_arith = "on";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~33 .shared_arith = "on";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~37 .shared_arith = "on";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~41 .shared_arith = "on";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout(\Add0~47 ));
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~45 .shared_arith = "on";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(\Add0~47 ),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout(\Add0~51 ));
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~49 .shared_arith = "on";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(\Add0~51 ),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout(\Add0~55 ));
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~53 .shared_arith = "on";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(\Add0~55 ),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout(\Add0~59 ));
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~57 .shared_arith = "on";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe162),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(\Add0~59 ),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout(\Add0~63 ));
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~61 .shared_arith = "on";

arriav_lcell_comb \Add0~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe171),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(\Add0~63 ),
	.combout(),
	.sumout(\Add0~65_sumout ),
	.cout(\Add0~66 ),
	.shareout(\Add0~67 ));
defparam \Add0~65 .extended_lut = "off";
defparam \Add0~65 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~65 .shared_arith = "on";

arriav_lcell_comb \Add0~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe181),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~66 ),
	.sharein(\Add0~67 ),
	.combout(),
	.sumout(\Add0~69_sumout ),
	.cout(),
	.shareout());
defparam \Add0~69 .extended_lut = "off";
defparam \Add0~69 .lut_mask = 64'h000000000000FF00;
defparam \Add0~69 .shared_arith = "on";

arriav_lcell_comb \xordvalue~0 (
	.dataa(!dffe161),
	.datab(!pipeline_dffe_17),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

endmodule

module nco_test_lpm_add_sub_34 (
	a_0,
	xordvalue_0,
	a_1,
	a_2,
	a_3,
	a_4,
	a_5,
	a_6,
	a_7,
	a_8,
	a_9,
	a_10,
	a_11,
	a_12,
	a_13,
	a_14,
	a_15,
	a_16,
	a_17,
	dffe1,
	dffe2,
	dffe3,
	dffe4,
	dffe5,
	dffe6,
	dffe7,
	dffe8,
	dffe9,
	dffe10,
	dffe11,
	dffe12,
	dffe13,
	dffe14,
	dffe15,
	dffe16,
	dffe17,
	dffe18,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_0;
input 	xordvalue_0;
input 	a_1;
input 	a_2;
input 	a_3;
input 	a_4;
input 	a_5;
input 	a_6;
input 	a_7;
input 	a_8;
input 	a_9;
input 	a_10;
input 	a_11;
input 	a_12;
input 	a_13;
input 	a_14;
input 	a_15;
input 	a_16;
input 	a_17;
output 	dffe1;
output 	dffe2;
output 	dffe3;
output 	dffe4;
output 	dffe5;
output 	dffe6;
output 	dffe7;
output 	dffe8;
output 	dffe9;
output 	dffe10;
output 	dffe11;
output 	dffe12;
output 	dffe13;
output 	dffe14;
output 	dffe15;
output 	dffe16;
output 	dffe17;
output 	dffe18;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_add_sub_jdg_15 auto_generated(
	.a_0(a_0),
	.xordvalue_0(xordvalue_0),
	.a_1(a_1),
	.a_2(a_2),
	.a_3(a_3),
	.a_4(a_4),
	.a_5(a_5),
	.a_6(a_6),
	.a_7(a_7),
	.a_8(a_8),
	.a_9(a_9),
	.a_10(a_10),
	.a_11(a_11),
	.a_12(a_12),
	.a_13(a_13),
	.a_14(a_14),
	.a_15(a_15),
	.a_16(a_16),
	.a_17(a_17),
	.dffe19(dffe1),
	.dffe21(dffe2),
	.dffe31(dffe3),
	.dffe41(dffe4),
	.dffe51(dffe5),
	.dffe61(dffe6),
	.dffe71(dffe7),
	.dffe81(dffe8),
	.dffe91(dffe9),
	.dffe101(dffe10),
	.dffe111(dffe11),
	.dffe121(dffe12),
	.dffe131(dffe13),
	.dffe141(dffe14),
	.dffe151(dffe15),
	.dffe161(dffe16),
	.dffe171(dffe17),
	.dffe181(dffe18),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module nco_test_add_sub_jdg_15 (
	a_0,
	xordvalue_0,
	a_1,
	a_2,
	a_3,
	a_4,
	a_5,
	a_6,
	a_7,
	a_8,
	a_9,
	a_10,
	a_11,
	a_12,
	a_13,
	a_14,
	a_15,
	a_16,
	a_17,
	dffe19,
	dffe21,
	dffe31,
	dffe41,
	dffe51,
	dffe61,
	dffe71,
	dffe81,
	dffe91,
	dffe101,
	dffe111,
	dffe121,
	dffe131,
	dffe141,
	dffe151,
	dffe161,
	dffe171,
	dffe181,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_0;
input 	xordvalue_0;
input 	a_1;
input 	a_2;
input 	a_3;
input 	a_4;
input 	a_5;
input 	a_6;
input 	a_7;
input 	a_8;
input 	a_9;
input 	a_10;
input 	a_11;
input 	a_12;
input 	a_13;
input 	a_14;
input 	a_15;
input 	a_16;
input 	a_17;
output 	dffe19;
output 	dffe21;
output 	dffe31;
output 	dffe41;
output 	dffe51;
output 	dffe61;
output 	dffe71;
output 	dffe81;
output 	dffe91;
output 	dffe101;
output 	dffe111;
output 	dffe121;
output 	dffe131;
output 	dffe141;
output 	dffe151;
output 	dffe161;
output 	dffe171;
output 	dffe181;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~sumout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~sumout ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~sumout ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~sumout ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~sumout ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~sumout ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~sumout ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~sumout ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~sumout ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~sumout ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~sumout ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~sumout ;
wire \add_sub_cella[11]~COUT ;
wire \add_sub_cella[12]~sumout ;
wire \add_sub_cella[12]~COUT ;
wire \add_sub_cella[13]~sumout ;
wire \add_sub_cella[13]~COUT ;
wire \add_sub_cella[14]~sumout ;
wire \add_sub_cella[14]~COUT ;
wire \add_sub_cella[15]~sumout ;
wire \add_sub_cella[15]~COUT ;
wire \add_sub_cella[16]~sumout ;
wire \add_sub_cella[16]~COUT ;
wire \add_sub_cella[17]~sumout ;


dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe19),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

dffeas dffe13(
	.clk(clock),
	.d(\add_sub_cella[12]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe131),
	.prn(vcc));
defparam dffe13.is_wysiwyg = "true";
defparam dffe13.power_up = "low";

dffeas dffe14(
	.clk(clock),
	.d(\add_sub_cella[13]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe141),
	.prn(vcc));
defparam dffe14.is_wysiwyg = "true";
defparam dffe14.power_up = "low";

dffeas dffe15(
	.clk(clock),
	.d(\add_sub_cella[14]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe151),
	.prn(vcc));
defparam dffe15.is_wysiwyg = "true";
defparam dffe15.power_up = "low";

dffeas dffe16(
	.clk(clock),
	.d(\add_sub_cella[15]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe161),
	.prn(vcc));
defparam dffe16.is_wysiwyg = "true";
defparam dffe16.power_up = "low";

dffeas dffe17(
	.clk(clock),
	.d(\add_sub_cella[16]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe171),
	.prn(vcc));
defparam dffe17.is_wysiwyg = "true";
defparam dffe17.power_up = "low";

dffeas dffe18(
	.clk(clock),
	.d(\add_sub_cella[17]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe181),
	.prn(vcc));
defparam dffe18.is_wysiwyg = "true";
defparam dffe18.power_up = "low";

arriav_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(\add_sub_cella[11]~COUT ),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[12] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[11]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[12]~sumout ),
	.cout(\add_sub_cella[12]~COUT ),
	.shareout());
defparam \add_sub_cella[12] .extended_lut = "off";
defparam \add_sub_cella[12] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[12] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[13] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[12]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[13]~sumout ),
	.cout(\add_sub_cella[13]~COUT ),
	.shareout());
defparam \add_sub_cella[13] .extended_lut = "off";
defparam \add_sub_cella[13] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[13] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[14] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[13]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[14]~sumout ),
	.cout(\add_sub_cella[14]~COUT ),
	.shareout());
defparam \add_sub_cella[14] .extended_lut = "off";
defparam \add_sub_cella[14] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[14] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[15] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[14]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[15]~sumout ),
	.cout(\add_sub_cella[15]~COUT ),
	.shareout());
defparam \add_sub_cella[15] .extended_lut = "off";
defparam \add_sub_cella[15] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[15] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[16] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_16),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[15]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[16]~sumout ),
	.cout(\add_sub_cella[16]~COUT ),
	.shareout());
defparam \add_sub_cella[16] .extended_lut = "off";
defparam \add_sub_cella[16] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[16] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[17] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_17),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[16]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[17]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[17] .extended_lut = "off";
defparam \add_sub_cella[17] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[17] .shared_arith = "off";

endmodule

module nco_test_cordic_sxor_1p_lpm_16 (
	sin_o_0,
	dffe18,
	dffe17,
	dffe16,
	pipeline_dffe_17,
	dffe161,
	dffe181,
	dffe15,
	pipeline_dffe_16,
	dffe171,
	dffe14,
	pipeline_dffe_15,
	dffe162,
	dffe13,
	pipeline_dffe_14,
	dffe151,
	dffe12,
	pipeline_dffe_13,
	dffe141,
	dffe11,
	pipeline_dffe_12,
	dffe131,
	dffe10,
	pipeline_dffe_11,
	dffe121,
	dffe9,
	pipeline_dffe_10,
	dffe111,
	dffe8,
	pipeline_dffe_9,
	dffe101,
	dffe7,
	pipeline_dffe_8,
	dffe91,
	dffe6,
	pipeline_dffe_7,
	dffe4,
	dffe5,
	dffe81,
	pipeline_dffe_6,
	dffe71,
	dffe1,
	pipeline_dffe_5,
	dffe2,
	dffe3,
	dffe61,
	pipeline_dffe_4,
	dffe51,
	pipeline_dffe_3,
	dffe31,
	dffe41,
	pipeline_dffe_2,
	dffe19,
	dffe21,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	sin_o_0;
output 	dffe18;
output 	dffe17;
input 	dffe16;
input 	pipeline_dffe_17;
output 	dffe161;
input 	dffe181;
output 	dffe15;
input 	pipeline_dffe_16;
input 	dffe171;
output 	dffe14;
input 	pipeline_dffe_15;
input 	dffe162;
output 	dffe13;
input 	pipeline_dffe_14;
input 	dffe151;
output 	dffe12;
input 	pipeline_dffe_13;
input 	dffe141;
output 	dffe11;
input 	pipeline_dffe_12;
input 	dffe131;
output 	dffe10;
input 	pipeline_dffe_11;
input 	dffe121;
output 	dffe9;
input 	pipeline_dffe_10;
input 	dffe111;
output 	dffe8;
input 	pipeline_dffe_9;
input 	dffe101;
output 	dffe7;
input 	pipeline_dffe_8;
input 	dffe91;
output 	dffe6;
input 	pipeline_dffe_7;
output 	dffe4;
output 	dffe5;
input 	dffe81;
input 	pipeline_dffe_6;
input 	dffe71;
output 	dffe1;
input 	pipeline_dffe_5;
output 	dffe2;
output 	dffe3;
input 	dffe61;
input 	pipeline_dffe_4;
input 	dffe51;
input 	pipeline_dffe_3;
input 	dffe31;
input 	dffe41;
input 	pipeline_dffe_2;
input 	dffe19;
input 	dffe21;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[17]~q ;
wire \xordvalue[15]~q ;
wire \Add0~1_sumout ;
wire \a[16]~q ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \a[15]~q ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \a[14]~q ;
wire \xordvalue[14]~q ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \a[13]~q ;
wire \xordvalue[13]~q ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \a[12]~q ;
wire \xordvalue[12]~q ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \a[11]~q ;
wire \xordvalue[11]~q ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \a[10]~q ;
wire \xordvalue[10]~q ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \a[9]~q ;
wire \xordvalue[9]~q ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \a[8]~q ;
wire \xordvalue[8]~q ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \a[7]~q ;
wire \xordvalue[7]~q ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \a[6]~q ;
wire \xordvalue[6]~q ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \a[5]~q ;
wire \xordvalue[5]~q ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~51 ;
wire \a[4]~q ;
wire \xordvalue[4]~q ;
wire \a[3]~q ;
wire \xordvalue[3]~q ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~55 ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~59 ;
wire \a[2]~q ;
wire \xordvalue[2]~q ;
wire \a[0]~q ;
wire \xordvalue[0]~q ;
wire \a[1]~q ;
wire \xordvalue[1]~q ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~63 ;
wire \Add0~65_sumout ;
wire \Add0~66 ;
wire \Add0~67 ;
wire \Add0~69_sumout ;
wire \Add0~70 ;
wire \Add0~71 ;
wire \xordvalue~0_combout ;
wire \xordvalue~1_combout ;
wire \xordvalue~2_combout ;
wire \xordvalue~3_combout ;
wire \xordvalue~4_combout ;
wire \xordvalue~5_combout ;
wire \xordvalue~6_combout ;
wire \xordvalue~7_combout ;
wire \xordvalue~8_combout ;
wire \xordvalue~9_combout ;
wire \xordvalue~10_combout ;
wire \xordvalue~11_combout ;
wire \xordvalue~12_combout ;
wire \xordvalue~13_combout ;
wire \xordvalue~14_combout ;
wire \xordvalue~15_combout ;


nco_test_lpm_add_sub_35 u0(
	.a_17(\a[17]~q ),
	.xordvalue_15(\xordvalue[15]~q ),
	.a_16(\a[16]~q ),
	.a_15(\a[15]~q ),
	.a_14(\a[14]~q ),
	.xordvalue_14(\xordvalue[14]~q ),
	.a_13(\a[13]~q ),
	.xordvalue_13(\xordvalue[13]~q ),
	.a_12(\a[12]~q ),
	.xordvalue_12(\xordvalue[12]~q ),
	.a_11(\a[11]~q ),
	.xordvalue_11(\xordvalue[11]~q ),
	.a_10(\a[10]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.a_9(\a[9]~q ),
	.xordvalue_9(\xordvalue[9]~q ),
	.a_8(\a[8]~q ),
	.xordvalue_8(\xordvalue[8]~q ),
	.a_7(\a[7]~q ),
	.xordvalue_7(\xordvalue[7]~q ),
	.a_6(\a[6]~q ),
	.xordvalue_6(\xordvalue[6]~q ),
	.a_5(\a[5]~q ),
	.xordvalue_5(\xordvalue[5]~q ),
	.a_4(\a[4]~q ),
	.xordvalue_4(\xordvalue[4]~q ),
	.a_3(\a[3]~q ),
	.xordvalue_3(\xordvalue[3]~q ),
	.a_2(\a[2]~q ),
	.xordvalue_2(\xordvalue[2]~q ),
	.a_0(\a[0]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_1(\a[1]~q ),
	.xordvalue_1(\xordvalue[1]~q ),
	.dffe18(dffe18),
	.dffe17(dffe17),
	.dffe16(dffe161),
	.dffe15(dffe15),
	.dffe14(dffe14),
	.dffe13(dffe13),
	.dffe12(dffe12),
	.dffe11(dffe11),
	.dffe10(dffe10),
	.dffe9(dffe9),
	.dffe8(dffe8),
	.dffe7(dffe7),
	.dffe6(dffe6),
	.dffe4(dffe4),
	.dffe5(dffe5),
	.dffe1(dffe1),
	.dffe2(dffe2),
	.dffe3(dffe3),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[17] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[17]~q ),
	.prn(vcc));
defparam \a[17] .is_wysiwyg = "true";
defparam \a[17] .power_up = "low";

dffeas \xordvalue[15] (
	.clk(clk),
	.d(\xordvalue~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[15]~q ),
	.prn(vcc));
defparam \xordvalue[15] .is_wysiwyg = "true";
defparam \xordvalue[15] .power_up = "low";

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe181),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "on";

dffeas \a[16] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[16]~q ),
	.prn(vcc));
defparam \a[16] .is_wysiwyg = "true";
defparam \a[16] .power_up = "low";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe171),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~5 .shared_arith = "on";

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe162),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~9 .shared_arith = "on";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

dffeas \xordvalue[14] (
	.clk(clk),
	.d(\xordvalue~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[14]~q ),
	.prn(vcc));
defparam \xordvalue[14] .is_wysiwyg = "true";
defparam \xordvalue[14] .power_up = "low";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~13 .shared_arith = "on";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

dffeas \xordvalue[13] (
	.clk(clk),
	.d(\xordvalue~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[13]~q ),
	.prn(vcc));
defparam \xordvalue[13] .is_wysiwyg = "true";
defparam \xordvalue[13] .power_up = "low";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~17 .shared_arith = "on";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

dffeas \xordvalue[12] (
	.clk(clk),
	.d(\xordvalue~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[12]~q ),
	.prn(vcc));
defparam \xordvalue[12] .is_wysiwyg = "true";
defparam \xordvalue[12] .power_up = "low";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "on";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \xordvalue[11] (
	.clk(clk),
	.d(\xordvalue~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[11]~q ),
	.prn(vcc));
defparam \xordvalue[11] .is_wysiwyg = "true";
defparam \xordvalue[11] .power_up = "low";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~25 .shared_arith = "on";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(\xordvalue~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~29 .shared_arith = "on";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \xordvalue[9] (
	.clk(clk),
	.d(\xordvalue~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[9]~q ),
	.prn(vcc));
defparam \xordvalue[9] .is_wysiwyg = "true";
defparam \xordvalue[9] .power_up = "low";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~33 .shared_arith = "on";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \xordvalue[8] (
	.clk(clk),
	.d(\xordvalue~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[8]~q ),
	.prn(vcc));
defparam \xordvalue[8] .is_wysiwyg = "true";
defparam \xordvalue[8] .power_up = "low";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~37 .shared_arith = "on";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \xordvalue[7] (
	.clk(clk),
	.d(\xordvalue~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[7]~q ),
	.prn(vcc));
defparam \xordvalue[7] .is_wysiwyg = "true";
defparam \xordvalue[7] .power_up = "low";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(\Add0~47 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~41 .shared_arith = "on";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \xordvalue[6] (
	.clk(clk),
	.d(\xordvalue~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[6]~q ),
	.prn(vcc));
defparam \xordvalue[6] .is_wysiwyg = "true";
defparam \xordvalue[6] .power_up = "low";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(\Add0~51 ),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout(\Add0~47 ));
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~45 .shared_arith = "on";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \xordvalue[5] (
	.clk(clk),
	.d(\xordvalue~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[5]~q ),
	.prn(vcc));
defparam \xordvalue[5] .is_wysiwyg = "true";
defparam \xordvalue[5] .power_up = "low";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(\Add0~55 ),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout(\Add0~51 ));
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~49 .shared_arith = "on";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \xordvalue[4] (
	.clk(clk),
	.d(\xordvalue~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[4]~q ),
	.prn(vcc));
defparam \xordvalue[4] .is_wysiwyg = "true";
defparam \xordvalue[4] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \xordvalue[3] (
	.clk(clk),
	.d(\xordvalue~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[3]~q ),
	.prn(vcc));
defparam \xordvalue[3] .is_wysiwyg = "true";
defparam \xordvalue[3] .power_up = "low";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(\Add0~59 ),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout(\Add0~55 ));
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~53 .shared_arith = "on";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(\Add0~63 ),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout(\Add0~59 ));
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~57 .shared_arith = "on";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \xordvalue[2] (
	.clk(clk),
	.d(\xordvalue~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[2]~q ),
	.prn(vcc));
defparam \xordvalue[2] .is_wysiwyg = "true";
defparam \xordvalue[2] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(\xordvalue~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \xordvalue[1] (
	.clk(clk),
	.d(\xordvalue~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[1]~q ),
	.prn(vcc));
defparam \xordvalue[1] .is_wysiwyg = "true";
defparam \xordvalue[1] .power_up = "low";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~70 ),
	.sharein(\Add0~71 ),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout(\Add0~63 ));
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~61 .shared_arith = "on";

arriav_lcell_comb \Add0~65 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!dffe19),
	.datad(!dffe16),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~65_sumout ),
	.cout(\Add0~66 ),
	.shareout(\Add0~67 ));
defparam \Add0~65 .extended_lut = "off";
defparam \Add0~65 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add0~65 .shared_arith = "on";

arriav_lcell_comb \Add0~69 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~66 ),
	.sharein(\Add0~67 ),
	.combout(),
	.sumout(\Add0~69_sumout ),
	.cout(\Add0~70 ),
	.shareout(\Add0~71 ));
defparam \Add0~69 .extended_lut = "off";
defparam \Add0~69 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~69 .shared_arith = "on";

arriav_lcell_comb \xordvalue~0 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_17),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~0_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~0 .extended_lut = "off";
defparam \xordvalue~0 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~0 .shared_arith = "off";

arriav_lcell_comb \xordvalue~1 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_16),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~1_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~1 .extended_lut = "off";
defparam \xordvalue~1 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~1 .shared_arith = "off";

arriav_lcell_comb \xordvalue~2 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_15),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~2_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~2 .extended_lut = "off";
defparam \xordvalue~2 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~2 .shared_arith = "off";

arriav_lcell_comb \xordvalue~3 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_14),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~3_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~3 .extended_lut = "off";
defparam \xordvalue~3 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~3 .shared_arith = "off";

arriav_lcell_comb \xordvalue~4 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_13),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~4_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~4 .extended_lut = "off";
defparam \xordvalue~4 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~4 .shared_arith = "off";

arriav_lcell_comb \xordvalue~5 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_12),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~5_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~5 .extended_lut = "off";
defparam \xordvalue~5 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~5 .shared_arith = "off";

arriav_lcell_comb \xordvalue~6 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_11),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~6_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~6 .extended_lut = "off";
defparam \xordvalue~6 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~6 .shared_arith = "off";

arriav_lcell_comb \xordvalue~7 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_10),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~7_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~7 .extended_lut = "off";
defparam \xordvalue~7 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~7 .shared_arith = "off";

arriav_lcell_comb \xordvalue~8 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_9),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~8_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~8 .extended_lut = "off";
defparam \xordvalue~8 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~8 .shared_arith = "off";

arriav_lcell_comb \xordvalue~9 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_8),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~9_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~9 .extended_lut = "off";
defparam \xordvalue~9 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~9 .shared_arith = "off";

arriav_lcell_comb \xordvalue~10 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_7),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~10_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~10 .extended_lut = "off";
defparam \xordvalue~10 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~10 .shared_arith = "off";

arriav_lcell_comb \xordvalue~11 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_6),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~11_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~11 .extended_lut = "off";
defparam \xordvalue~11 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~11 .shared_arith = "off";

arriav_lcell_comb \xordvalue~12 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_5),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~12_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~12 .extended_lut = "off";
defparam \xordvalue~12 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~12 .shared_arith = "off";

arriav_lcell_comb \xordvalue~13 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_4),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~13_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~13 .extended_lut = "off";
defparam \xordvalue~13 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~13 .shared_arith = "off";

arriav_lcell_comb \xordvalue~14 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_2),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~14_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~14 .extended_lut = "off";
defparam \xordvalue~14 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~14 .shared_arith = "off";

arriav_lcell_comb \xordvalue~15 (
	.dataa(!dffe16),
	.datab(!pipeline_dffe_3),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(\xordvalue~15_combout ),
	.sumout(),
	.cout(),
	.shareout());
defparam \xordvalue~15 .extended_lut = "off";
defparam \xordvalue~15 .lut_mask = 64'h6666666666666666;
defparam \xordvalue~15 .shared_arith = "off";

endmodule

module nco_test_lpm_add_sub_35 (
	a_17,
	xordvalue_15,
	a_16,
	a_15,
	a_14,
	xordvalue_14,
	a_13,
	xordvalue_13,
	a_12,
	xordvalue_12,
	a_11,
	xordvalue_11,
	a_10,
	xordvalue_10,
	a_9,
	xordvalue_9,
	a_8,
	xordvalue_8,
	a_7,
	xordvalue_7,
	a_6,
	xordvalue_6,
	a_5,
	xordvalue_5,
	a_4,
	xordvalue_4,
	a_3,
	xordvalue_3,
	a_2,
	xordvalue_2,
	a_0,
	xordvalue_0,
	a_1,
	xordvalue_1,
	dffe18,
	dffe17,
	dffe16,
	dffe15,
	dffe14,
	dffe13,
	dffe12,
	dffe11,
	dffe10,
	dffe9,
	dffe8,
	dffe7,
	dffe6,
	dffe4,
	dffe5,
	dffe1,
	dffe2,
	dffe3,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_15;
input 	a_16;
input 	a_15;
input 	a_14;
input 	xordvalue_14;
input 	a_13;
input 	xordvalue_13;
input 	a_12;
input 	xordvalue_12;
input 	a_11;
input 	xordvalue_11;
input 	a_10;
input 	xordvalue_10;
input 	a_9;
input 	xordvalue_9;
input 	a_8;
input 	xordvalue_8;
input 	a_7;
input 	xordvalue_7;
input 	a_6;
input 	xordvalue_6;
input 	a_5;
input 	xordvalue_5;
input 	a_4;
input 	xordvalue_4;
input 	a_3;
input 	xordvalue_3;
input 	a_2;
input 	xordvalue_2;
input 	a_0;
input 	xordvalue_0;
input 	a_1;
input 	xordvalue_1;
output 	dffe18;
output 	dffe17;
output 	dffe16;
output 	dffe15;
output 	dffe14;
output 	dffe13;
output 	dffe12;
output 	dffe11;
output 	dffe10;
output 	dffe9;
output 	dffe8;
output 	dffe7;
output 	dffe6;
output 	dffe4;
output 	dffe5;
output 	dffe1;
output 	dffe2;
output 	dffe3;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_add_sub_jdg_16 auto_generated(
	.a_17(a_17),
	.xordvalue_15(xordvalue_15),
	.a_16(a_16),
	.a_15(a_15),
	.a_14(a_14),
	.xordvalue_14(xordvalue_14),
	.a_13(a_13),
	.xordvalue_13(xordvalue_13),
	.a_12(a_12),
	.xordvalue_12(xordvalue_12),
	.a_11(a_11),
	.xordvalue_11(xordvalue_11),
	.a_10(a_10),
	.xordvalue_10(xordvalue_10),
	.a_9(a_9),
	.xordvalue_9(xordvalue_9),
	.a_8(a_8),
	.xordvalue_8(xordvalue_8),
	.a_7(a_7),
	.xordvalue_7(xordvalue_7),
	.a_6(a_6),
	.xordvalue_6(xordvalue_6),
	.a_5(a_5),
	.xordvalue_5(xordvalue_5),
	.a_4(a_4),
	.xordvalue_4(xordvalue_4),
	.a_3(a_3),
	.xordvalue_3(xordvalue_3),
	.a_2(a_2),
	.xordvalue_2(xordvalue_2),
	.a_0(a_0),
	.xordvalue_0(xordvalue_0),
	.a_1(a_1),
	.xordvalue_1(xordvalue_1),
	.dffe181(dffe18),
	.dffe171(dffe17),
	.dffe161(dffe16),
	.dffe151(dffe15),
	.dffe141(dffe14),
	.dffe131(dffe13),
	.dffe121(dffe12),
	.dffe111(dffe11),
	.dffe101(dffe10),
	.dffe91(dffe9),
	.dffe81(dffe8),
	.dffe71(dffe7),
	.dffe61(dffe6),
	.dffe41(dffe4),
	.dffe51(dffe5),
	.dffe19(dffe1),
	.dffe21(dffe2),
	.dffe31(dffe3),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module nco_test_add_sub_jdg_16 (
	a_17,
	xordvalue_15,
	a_16,
	a_15,
	a_14,
	xordvalue_14,
	a_13,
	xordvalue_13,
	a_12,
	xordvalue_12,
	a_11,
	xordvalue_11,
	a_10,
	xordvalue_10,
	a_9,
	xordvalue_9,
	a_8,
	xordvalue_8,
	a_7,
	xordvalue_7,
	a_6,
	xordvalue_6,
	a_5,
	xordvalue_5,
	a_4,
	xordvalue_4,
	a_3,
	xordvalue_3,
	a_2,
	xordvalue_2,
	a_0,
	xordvalue_0,
	a_1,
	xordvalue_1,
	dffe181,
	dffe171,
	dffe161,
	dffe151,
	dffe141,
	dffe131,
	dffe121,
	dffe111,
	dffe101,
	dffe91,
	dffe81,
	dffe71,
	dffe61,
	dffe41,
	dffe51,
	dffe19,
	dffe21,
	dffe31,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_17;
input 	xordvalue_15;
input 	a_16;
input 	a_15;
input 	a_14;
input 	xordvalue_14;
input 	a_13;
input 	xordvalue_13;
input 	a_12;
input 	xordvalue_12;
input 	a_11;
input 	xordvalue_11;
input 	a_10;
input 	xordvalue_10;
input 	a_9;
input 	xordvalue_9;
input 	a_8;
input 	xordvalue_8;
input 	a_7;
input 	xordvalue_7;
input 	a_6;
input 	xordvalue_6;
input 	a_5;
input 	xordvalue_5;
input 	a_4;
input 	xordvalue_4;
input 	a_3;
input 	xordvalue_3;
input 	a_2;
input 	xordvalue_2;
input 	a_0;
input 	xordvalue_0;
input 	a_1;
input 	xordvalue_1;
output 	dffe181;
output 	dffe171;
output 	dffe161;
output 	dffe151;
output 	dffe141;
output 	dffe131;
output 	dffe121;
output 	dffe111;
output 	dffe101;
output 	dffe91;
output 	dffe81;
output 	dffe71;
output 	dffe61;
output 	dffe41;
output 	dffe51;
output 	dffe19;
output 	dffe21;
output 	dffe31;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~COUT ;
wire \add_sub_cella[12]~COUT ;
wire \add_sub_cella[13]~COUT ;
wire \add_sub_cella[14]~COUT ;
wire \add_sub_cella[15]~COUT ;
wire \add_sub_cella[16]~COUT ;
wire \add_sub_cella[17]~sumout ;
wire \add_sub_cella[16]~sumout ;
wire \add_sub_cella[15]~sumout ;
wire \add_sub_cella[14]~sumout ;
wire \add_sub_cella[13]~sumout ;
wire \add_sub_cella[12]~sumout ;
wire \add_sub_cella[11]~sumout ;
wire \add_sub_cella[10]~sumout ;
wire \add_sub_cella[9]~sumout ;
wire \add_sub_cella[8]~sumout ;
wire \add_sub_cella[7]~sumout ;
wire \add_sub_cella[6]~sumout ;
wire \add_sub_cella[5]~sumout ;
wire \add_sub_cella[3]~sumout ;
wire \add_sub_cella[4]~sumout ;
wire \add_sub_cella[0]~sumout ;
wire \add_sub_cella[1]~sumout ;
wire \add_sub_cella[2]~sumout ;


dffeas dffe18(
	.clk(clock),
	.d(\add_sub_cella[17]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe181),
	.prn(vcc));
defparam dffe18.is_wysiwyg = "true";
defparam dffe18.power_up = "low";

dffeas dffe17(
	.clk(clock),
	.d(\add_sub_cella[16]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe171),
	.prn(vcc));
defparam dffe17.is_wysiwyg = "true";
defparam dffe17.power_up = "low";

dffeas dffe16(
	.clk(clock),
	.d(\add_sub_cella[15]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe161),
	.prn(vcc));
defparam dffe16.is_wysiwyg = "true";
defparam dffe16.power_up = "low";

dffeas dffe15(
	.clk(clock),
	.d(\add_sub_cella[14]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe151),
	.prn(vcc));
defparam dffe15.is_wysiwyg = "true";
defparam dffe15.power_up = "low";

dffeas dffe14(
	.clk(clock),
	.d(\add_sub_cella[13]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe141),
	.prn(vcc));
defparam dffe14.is_wysiwyg = "true";
defparam dffe14.power_up = "low";

dffeas dffe13(
	.clk(clock),
	.d(\add_sub_cella[12]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe131),
	.prn(vcc));
defparam dffe13.is_wysiwyg = "true";
defparam dffe13.power_up = "low";

dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe19),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

arriav_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_1),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_2),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_3),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_4),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_5),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_6),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_7),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_8),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_9),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_11),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(\add_sub_cella[11]~COUT ),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[12] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_12),
	.datag(gnd),
	.cin(\add_sub_cella[11]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[12]~sumout ),
	.cout(\add_sub_cella[12]~COUT ),
	.shareout());
defparam \add_sub_cella[12] .extended_lut = "off";
defparam \add_sub_cella[12] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[12] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[13] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_13),
	.datag(gnd),
	.cin(\add_sub_cella[12]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[13]~sumout ),
	.cout(\add_sub_cella[13]~COUT ),
	.shareout());
defparam \add_sub_cella[13] .extended_lut = "off";
defparam \add_sub_cella[13] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[13] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[14] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_14),
	.datag(gnd),
	.cin(\add_sub_cella[13]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[14]~sumout ),
	.cout(\add_sub_cella[14]~COUT ),
	.shareout());
defparam \add_sub_cella[14] .extended_lut = "off";
defparam \add_sub_cella[14] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[14] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[15] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_15),
	.datag(gnd),
	.cin(\add_sub_cella[14]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[15]~sumout ),
	.cout(\add_sub_cella[15]~COUT ),
	.shareout());
defparam \add_sub_cella[15] .extended_lut = "off";
defparam \add_sub_cella[15] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[15] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[16] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_16),
	.datae(gnd),
	.dataf(!xordvalue_15),
	.datag(gnd),
	.cin(\add_sub_cella[15]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[16]~sumout ),
	.cout(\add_sub_cella[16]~COUT ),
	.shareout());
defparam \add_sub_cella[16] .extended_lut = "off";
defparam \add_sub_cella[16] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[16] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[17] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_17),
	.datae(gnd),
	.dataf(!xordvalue_15),
	.datag(gnd),
	.cin(\add_sub_cella[16]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[17]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[17] .extended_lut = "off";
defparam \add_sub_cella[17] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[17] .shared_arith = "off";

endmodule

module nco_test_cordic_zxor_1p_lpm (
	sin_o_0,
	dffe16,
	dffe15,
	dffe14,
	dffe161,
	dffe13,
	dffe12,
	dffe151,
	dffe11,
	dffe141,
	dffe10,
	dffe131,
	dffe9,
	dffe121,
	dffe8,
	dffe111,
	dffe7,
	dffe101,
	dffe6,
	dffe91,
	dffe5,
	dffe81,
	dffe4,
	dffe71,
	dffe3,
	dffe61,
	dffe2,
	dffe51,
	dffe1,
	dffe41,
	dffe31,
	dffe21,
	dffe17,
	dffe162,
	dffe163,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	sin_o_0;
output 	dffe16;
output 	dffe15;
output 	dffe14;
input 	dffe161;
output 	dffe13;
output 	dffe12;
input 	dffe151;
output 	dffe11;
input 	dffe141;
output 	dffe10;
input 	dffe131;
output 	dffe9;
input 	dffe121;
output 	dffe8;
input 	dffe111;
output 	dffe7;
input 	dffe101;
output 	dffe6;
input 	dffe91;
output 	dffe5;
input 	dffe81;
output 	dffe4;
input 	dffe71;
output 	dffe3;
input 	dffe61;
output 	dffe2;
input 	dffe51;
output 	dffe1;
input 	dffe41;
input 	dffe31;
input 	dffe21;
input 	dffe17;
output 	dffe162;
input 	dffe163;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[15]~q ;
wire \xordvalue[0]~q ;
wire \Add0~1_sumout ;
wire \a[14]~q ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \a[13]~q ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \a[12]~q ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \a[11]~q ;
wire \xordvalue[11]~q ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \a[10]~q ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \a[9]~q ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \a[8]~q ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \a[7]~q ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \a[6]~q ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \a[5]~q ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \a[4]~q ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \a[3]~q ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~51 ;
wire \a[2]~q ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~55 ;
wire \a[1]~q ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~59 ;
wire \a[0]~q ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~63 ;


nco_test_lpm_add_sub_36 u0(
	.a_15(\a[15]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_14(\a[14]~q ),
	.a_13(\a[13]~q ),
	.a_12(\a[12]~q ),
	.a_11(\a[11]~q ),
	.xordvalue_11(\xordvalue[11]~q ),
	.a_10(\a[10]~q ),
	.a_9(\a[9]~q ),
	.a_8(\a[8]~q ),
	.a_7(\a[7]~q ),
	.a_6(\a[6]~q ),
	.a_5(\a[5]~q ),
	.a_4(\a[4]~q ),
	.a_3(\a[3]~q ),
	.a_2(\a[2]~q ),
	.a_1(\a[1]~q ),
	.a_0(\a[0]~q ),
	.dffe16(dffe16),
	.dffe15(dffe15),
	.dffe14(dffe14),
	.dffe13(dffe13),
	.dffe12(dffe12),
	.dffe11(dffe11),
	.dffe10(dffe10),
	.dffe9(dffe9),
	.dffe8(dffe8),
	.dffe7(dffe7),
	.dffe6(dffe6),
	.dffe5(dffe5),
	.dffe4(dffe4),
	.dffe3(dffe3),
	.dffe2(dffe2),
	.dffe1(dffe1),
	.dffe161(dffe162),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(dffe161),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "on";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~5 .shared_arith = "on";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~9 .shared_arith = "on";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~13 .shared_arith = "on";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \xordvalue[11] (
	.clk(clk),
	.d(dffe163),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[11]~q ),
	.prn(vcc));
defparam \xordvalue[11] .is_wysiwyg = "true";
defparam \xordvalue[11] .power_up = "low";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~17 .shared_arith = "on";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "on";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~25 .shared_arith = "on";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~29 .shared_arith = "on";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~33 .shared_arith = "on";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~37 .shared_arith = "on";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(\Add0~47 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~41 .shared_arith = "on";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(\Add0~51 ),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout(\Add0~47 ));
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~45 .shared_arith = "on";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(\Add0~55 ),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout(\Add0~51 ));
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~49 .shared_arith = "on";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(\Add0~59 ),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout(\Add0~55 ));
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~53 .shared_arith = "on";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(\Add0~63 ),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout(\Add0~59 ));
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~57 .shared_arith = "on";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!dffe17),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout(\Add0~63 ));
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add0~61 .shared_arith = "on";

endmodule

module nco_test_lpm_add_sub_36 (
	a_15,
	xordvalue_0,
	a_14,
	a_13,
	a_12,
	a_11,
	xordvalue_11,
	a_10,
	a_9,
	a_8,
	a_7,
	a_6,
	a_5,
	a_4,
	a_3,
	a_2,
	a_1,
	a_0,
	dffe16,
	dffe15,
	dffe14,
	dffe13,
	dffe12,
	dffe11,
	dffe10,
	dffe9,
	dffe8,
	dffe7,
	dffe6,
	dffe5,
	dffe4,
	dffe3,
	dffe2,
	dffe1,
	dffe161,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_15;
input 	xordvalue_0;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	xordvalue_11;
input 	a_10;
input 	a_9;
input 	a_8;
input 	a_7;
input 	a_6;
input 	a_5;
input 	a_4;
input 	a_3;
input 	a_2;
input 	a_1;
input 	a_0;
output 	dffe16;
output 	dffe15;
output 	dffe14;
output 	dffe13;
output 	dffe12;
output 	dffe11;
output 	dffe10;
output 	dffe9;
output 	dffe8;
output 	dffe7;
output 	dffe6;
output 	dffe5;
output 	dffe4;
output 	dffe3;
output 	dffe2;
output 	dffe1;
output 	dffe161;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_add_sub_hdg auto_generated(
	.a_15(a_15),
	.xordvalue_0(xordvalue_0),
	.a_14(a_14),
	.a_13(a_13),
	.a_12(a_12),
	.a_11(a_11),
	.xordvalue_11(xordvalue_11),
	.a_10(a_10),
	.a_9(a_9),
	.a_8(a_8),
	.a_7(a_7),
	.a_6(a_6),
	.a_5(a_5),
	.a_4(a_4),
	.a_3(a_3),
	.a_2(a_2),
	.a_1(a_1),
	.a_0(a_0),
	.dffe161(dffe16),
	.dffe151(dffe15),
	.dffe141(dffe14),
	.dffe131(dffe13),
	.dffe121(dffe12),
	.dffe111(dffe11),
	.dffe101(dffe10),
	.dffe91(dffe9),
	.dffe81(dffe8),
	.dffe71(dffe7),
	.dffe61(dffe6),
	.dffe51(dffe5),
	.dffe41(dffe4),
	.dffe31(dffe3),
	.dffe21(dffe2),
	.dffe17(dffe1),
	.dffe162(dffe161),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module nco_test_add_sub_hdg (
	a_15,
	xordvalue_0,
	a_14,
	a_13,
	a_12,
	a_11,
	xordvalue_11,
	a_10,
	a_9,
	a_8,
	a_7,
	a_6,
	a_5,
	a_4,
	a_3,
	a_2,
	a_1,
	a_0,
	dffe161,
	dffe151,
	dffe141,
	dffe131,
	dffe121,
	dffe111,
	dffe101,
	dffe91,
	dffe81,
	dffe71,
	dffe61,
	dffe51,
	dffe41,
	dffe31,
	dffe21,
	dffe17,
	dffe162,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_15;
input 	xordvalue_0;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	xordvalue_11;
input 	a_10;
input 	a_9;
input 	a_8;
input 	a_7;
input 	a_6;
input 	a_5;
input 	a_4;
input 	a_3;
input 	a_2;
input 	a_1;
input 	a_0;
output 	dffe161;
output 	dffe151;
output 	dffe141;
output 	dffe131;
output 	dffe121;
output 	dffe111;
output 	dffe101;
output 	dffe91;
output 	dffe81;
output 	dffe71;
output 	dffe61;
output 	dffe51;
output 	dffe41;
output 	dffe31;
output 	dffe21;
output 	dffe17;
output 	dffe162;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~COUT ;
wire \add_sub_cella[12]~COUT ;
wire \add_sub_cella[13]~COUT ;
wire \add_sub_cella[14]~COUT ;
wire \add_sub_cella[15]~sumout ;
wire \add_sub_cella[14]~sumout ;
wire \add_sub_cella[13]~sumout ;
wire \add_sub_cella[12]~sumout ;
wire \add_sub_cella[11]~sumout ;
wire \add_sub_cella[10]~sumout ;
wire \add_sub_cella[9]~sumout ;
wire \add_sub_cella[8]~sumout ;
wire \add_sub_cella[7]~sumout ;
wire \add_sub_cella[6]~sumout ;
wire \add_sub_cella[5]~sumout ;
wire \add_sub_cella[4]~sumout ;
wire \add_sub_cella[3]~sumout ;
wire \add_sub_cella[2]~sumout ;
wire \add_sub_cella[1]~sumout ;
wire \add_sub_cella[0]~sumout ;


dffeas dffe16(
	.clk(clock),
	.d(\add_sub_cella[15]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe161),
	.prn(vcc));
defparam dffe16.is_wysiwyg = "true";
defparam dffe16.power_up = "low";

dffeas dffe15(
	.clk(clock),
	.d(\add_sub_cella[14]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe151),
	.prn(vcc));
defparam dffe15.is_wysiwyg = "true";
defparam dffe15.power_up = "low";

dffeas dffe14(
	.clk(clock),
	.d(\add_sub_cella[13]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe141),
	.prn(vcc));
defparam dffe14.is_wysiwyg = "true";
defparam dffe14.power_up = "low";

dffeas dffe13(
	.clk(clock),
	.d(\add_sub_cella[12]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe131),
	.prn(vcc));
defparam dffe13.is_wysiwyg = "true";
defparam dffe13.power_up = "low";

dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe17),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

arriav_lcell_comb \dffe16~_wirecell (
	.dataa(!dffe161),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(dffe162),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffe16~_wirecell .extended_lut = "off";
defparam \dffe16~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dffe16~_wirecell .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_11),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_11),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_11),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_11),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(\add_sub_cella[11]~COUT ),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[12] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[11]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[12]~sumout ),
	.cout(\add_sub_cella[12]~COUT ),
	.shareout());
defparam \add_sub_cella[12] .extended_lut = "off";
defparam \add_sub_cella[12] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[12] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[13] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[12]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[13]~sumout ),
	.cout(\add_sub_cella[13]~COUT ),
	.shareout());
defparam \add_sub_cella[13] .extended_lut = "off";
defparam \add_sub_cella[13] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[13] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[14] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[13]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[14]~sumout ),
	.cout(\add_sub_cella[14]~COUT ),
	.shareout());
defparam \add_sub_cella[14] .extended_lut = "off";
defparam \add_sub_cella[14] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[14] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[15] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[14]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[15]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[15] .extended_lut = "off";
defparam \add_sub_cella[15] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[15] .shared_arith = "off";

endmodule

module nco_test_cordic_zxor_1p_lpm_1 (
	sin_o_0,
	dffe16,
	dffe15,
	dffe14,
	dffe161,
	dffe13,
	dffe12,
	dffe151,
	dffe11,
	dffe141,
	dffe10,
	dffe131,
	dffe9,
	dffe121,
	dffe8,
	dffe111,
	dffe7,
	dffe101,
	dffe6,
	dffe91,
	dffe5,
	dffe81,
	dffe4,
	dffe71,
	dffe3,
	dffe61,
	dffe2,
	dffe51,
	dffe1,
	dffe41,
	dffe31,
	dffe21,
	dffe17,
	dffe162,
	dffe163,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	sin_o_0;
output 	dffe16;
output 	dffe15;
output 	dffe14;
input 	dffe161;
output 	dffe13;
output 	dffe12;
input 	dffe151;
output 	dffe11;
input 	dffe141;
output 	dffe10;
input 	dffe131;
output 	dffe9;
input 	dffe121;
output 	dffe8;
input 	dffe111;
output 	dffe7;
input 	dffe101;
output 	dffe6;
input 	dffe91;
output 	dffe5;
input 	dffe81;
output 	dffe4;
input 	dffe71;
output 	dffe3;
input 	dffe61;
output 	dffe2;
input 	dffe51;
output 	dffe1;
input 	dffe41;
input 	dffe31;
input 	dffe21;
input 	dffe17;
input 	dffe162;
output 	dffe163;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[15]~q ;
wire \xordvalue[0]~q ;
wire \Add0~1_sumout ;
wire \a[14]~q ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \a[13]~q ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \a[12]~q ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \a[11]~q ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \a[10]~q ;
wire \xordvalue[10]~q ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \a[9]~q ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \a[8]~q ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \a[7]~q ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \a[6]~q ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \a[5]~q ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \a[4]~q ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \a[3]~q ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~51 ;
wire \a[2]~q ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~55 ;
wire \a[1]~q ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~59 ;
wire \a[0]~q ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~63 ;


nco_test_lpm_add_sub_37 u0(
	.a_15(\a[15]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_14(\a[14]~q ),
	.a_13(\a[13]~q ),
	.a_12(\a[12]~q ),
	.a_11(\a[11]~q ),
	.a_10(\a[10]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.a_9(\a[9]~q ),
	.a_8(\a[8]~q ),
	.a_7(\a[7]~q ),
	.a_6(\a[6]~q ),
	.a_5(\a[5]~q ),
	.a_4(\a[4]~q ),
	.a_3(\a[3]~q ),
	.a_2(\a[2]~q ),
	.a_1(\a[1]~q ),
	.a_0(\a[0]~q ),
	.dffe16(dffe16),
	.dffe15(dffe15),
	.dffe14(dffe14),
	.dffe13(dffe13),
	.dffe12(dffe12),
	.dffe11(dffe11),
	.dffe10(dffe10),
	.dffe9(dffe9),
	.dffe8(dffe8),
	.dffe7(dffe7),
	.dffe6(dffe6),
	.dffe5(dffe5),
	.dffe4(dffe4),
	.dffe3(dffe3),
	.dffe2(dffe2),
	.dffe1(dffe1),
	.dffe161(dffe163),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(dffe161),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "on";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~5 .shared_arith = "on";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~9 .shared_arith = "on";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~13 .shared_arith = "on";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~17 .shared_arith = "on";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(dffe162),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "on";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~25 .shared_arith = "on";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~29 .shared_arith = "on";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~33 .shared_arith = "on";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~37 .shared_arith = "on";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(\Add0~47 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~41 .shared_arith = "on";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(\Add0~51 ),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout(\Add0~47 ));
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~45 .shared_arith = "on";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(\Add0~55 ),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout(\Add0~51 ));
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~49 .shared_arith = "on";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(\Add0~59 ),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout(\Add0~55 ));
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~53 .shared_arith = "on";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(\Add0~63 ),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout(\Add0~59 ));
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~57 .shared_arith = "on";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!dffe17),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout(\Add0~63 ));
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add0~61 .shared_arith = "on";

endmodule

module nco_test_lpm_add_sub_37 (
	a_15,
	xordvalue_0,
	a_14,
	a_13,
	a_12,
	a_11,
	a_10,
	xordvalue_10,
	a_9,
	a_8,
	a_7,
	a_6,
	a_5,
	a_4,
	a_3,
	a_2,
	a_1,
	a_0,
	dffe16,
	dffe15,
	dffe14,
	dffe13,
	dffe12,
	dffe11,
	dffe10,
	dffe9,
	dffe8,
	dffe7,
	dffe6,
	dffe5,
	dffe4,
	dffe3,
	dffe2,
	dffe1,
	dffe161,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_15;
input 	xordvalue_0;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_10;
input 	xordvalue_10;
input 	a_9;
input 	a_8;
input 	a_7;
input 	a_6;
input 	a_5;
input 	a_4;
input 	a_3;
input 	a_2;
input 	a_1;
input 	a_0;
output 	dffe16;
output 	dffe15;
output 	dffe14;
output 	dffe13;
output 	dffe12;
output 	dffe11;
output 	dffe10;
output 	dffe9;
output 	dffe8;
output 	dffe7;
output 	dffe6;
output 	dffe5;
output 	dffe4;
output 	dffe3;
output 	dffe2;
output 	dffe1;
output 	dffe161;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_add_sub_hdg_1 auto_generated(
	.a_15(a_15),
	.xordvalue_0(xordvalue_0),
	.a_14(a_14),
	.a_13(a_13),
	.a_12(a_12),
	.a_11(a_11),
	.a_10(a_10),
	.xordvalue_10(xordvalue_10),
	.a_9(a_9),
	.a_8(a_8),
	.a_7(a_7),
	.a_6(a_6),
	.a_5(a_5),
	.a_4(a_4),
	.a_3(a_3),
	.a_2(a_2),
	.a_1(a_1),
	.a_0(a_0),
	.dffe161(dffe16),
	.dffe151(dffe15),
	.dffe141(dffe14),
	.dffe131(dffe13),
	.dffe121(dffe12),
	.dffe111(dffe11),
	.dffe101(dffe10),
	.dffe91(dffe9),
	.dffe81(dffe8),
	.dffe71(dffe7),
	.dffe61(dffe6),
	.dffe51(dffe5),
	.dffe41(dffe4),
	.dffe31(dffe3),
	.dffe21(dffe2),
	.dffe17(dffe1),
	.dffe162(dffe161),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module nco_test_add_sub_hdg_1 (
	a_15,
	xordvalue_0,
	a_14,
	a_13,
	a_12,
	a_11,
	a_10,
	xordvalue_10,
	a_9,
	a_8,
	a_7,
	a_6,
	a_5,
	a_4,
	a_3,
	a_2,
	a_1,
	a_0,
	dffe161,
	dffe151,
	dffe141,
	dffe131,
	dffe121,
	dffe111,
	dffe101,
	dffe91,
	dffe81,
	dffe71,
	dffe61,
	dffe51,
	dffe41,
	dffe31,
	dffe21,
	dffe17,
	dffe162,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_15;
input 	xordvalue_0;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_10;
input 	xordvalue_10;
input 	a_9;
input 	a_8;
input 	a_7;
input 	a_6;
input 	a_5;
input 	a_4;
input 	a_3;
input 	a_2;
input 	a_1;
input 	a_0;
output 	dffe161;
output 	dffe151;
output 	dffe141;
output 	dffe131;
output 	dffe121;
output 	dffe111;
output 	dffe101;
output 	dffe91;
output 	dffe81;
output 	dffe71;
output 	dffe61;
output 	dffe51;
output 	dffe41;
output 	dffe31;
output 	dffe21;
output 	dffe17;
output 	dffe162;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~COUT ;
wire \add_sub_cella[12]~COUT ;
wire \add_sub_cella[13]~COUT ;
wire \add_sub_cella[14]~COUT ;
wire \add_sub_cella[15]~sumout ;
wire \add_sub_cella[14]~sumout ;
wire \add_sub_cella[13]~sumout ;
wire \add_sub_cella[12]~sumout ;
wire \add_sub_cella[11]~sumout ;
wire \add_sub_cella[10]~sumout ;
wire \add_sub_cella[9]~sumout ;
wire \add_sub_cella[8]~sumout ;
wire \add_sub_cella[7]~sumout ;
wire \add_sub_cella[6]~sumout ;
wire \add_sub_cella[5]~sumout ;
wire \add_sub_cella[4]~sumout ;
wire \add_sub_cella[3]~sumout ;
wire \add_sub_cella[2]~sumout ;
wire \add_sub_cella[1]~sumout ;
wire \add_sub_cella[0]~sumout ;


dffeas dffe16(
	.clk(clock),
	.d(\add_sub_cella[15]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe161),
	.prn(vcc));
defparam dffe16.is_wysiwyg = "true";
defparam dffe16.power_up = "low";

dffeas dffe15(
	.clk(clock),
	.d(\add_sub_cella[14]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe151),
	.prn(vcc));
defparam dffe15.is_wysiwyg = "true";
defparam dffe15.power_up = "low";

dffeas dffe14(
	.clk(clock),
	.d(\add_sub_cella[13]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe141),
	.prn(vcc));
defparam dffe14.is_wysiwyg = "true";
defparam dffe14.power_up = "low";

dffeas dffe13(
	.clk(clock),
	.d(\add_sub_cella[12]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe131),
	.prn(vcc));
defparam dffe13.is_wysiwyg = "true";
defparam dffe13.power_up = "low";

dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe17),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

arriav_lcell_comb \dffe16~_wirecell (
	.dataa(!dffe161),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(dffe162),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffe16~_wirecell .extended_lut = "off";
defparam \dffe16~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dffe16~_wirecell .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(\add_sub_cella[11]~COUT ),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[12] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[11]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[12]~sumout ),
	.cout(\add_sub_cella[12]~COUT ),
	.shareout());
defparam \add_sub_cella[12] .extended_lut = "off";
defparam \add_sub_cella[12] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[12] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[13] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[12]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[13]~sumout ),
	.cout(\add_sub_cella[13]~COUT ),
	.shareout());
defparam \add_sub_cella[13] .extended_lut = "off";
defparam \add_sub_cella[13] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[13] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[14] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[13]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[14]~sumout ),
	.cout(\add_sub_cella[14]~COUT ),
	.shareout());
defparam \add_sub_cella[14] .extended_lut = "off";
defparam \add_sub_cella[14] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[14] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[15] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[14]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[15]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[15] .extended_lut = "off";
defparam \add_sub_cella[15] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[15] .shared_arith = "off";

endmodule

module nco_test_cordic_zxor_1p_lpm_2 (
	sin_o_0,
	dffe16,
	dffe15,
	dffe14,
	dffe161,
	dffe13,
	dffe12,
	dffe151,
	dffe11,
	dffe141,
	dffe10,
	dffe131,
	dffe9,
	dffe121,
	dffe8,
	dffe111,
	dffe7,
	dffe101,
	dffe6,
	dffe91,
	dffe5,
	dffe81,
	dffe4,
	dffe71,
	dffe3,
	dffe61,
	dffe2,
	dffe51,
	dffe1,
	dffe41,
	dffe31,
	dffe21,
	dffe17,
	dffe162,
	dffe163,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	sin_o_0;
output 	dffe16;
output 	dffe15;
output 	dffe14;
input 	dffe161;
output 	dffe13;
output 	dffe12;
input 	dffe151;
output 	dffe11;
input 	dffe141;
output 	dffe10;
input 	dffe131;
output 	dffe9;
input 	dffe121;
output 	dffe8;
input 	dffe111;
output 	dffe7;
input 	dffe101;
output 	dffe6;
input 	dffe91;
output 	dffe5;
input 	dffe81;
output 	dffe4;
input 	dffe71;
output 	dffe3;
input 	dffe61;
output 	dffe2;
input 	dffe51;
output 	dffe1;
input 	dffe41;
input 	dffe31;
input 	dffe21;
input 	dffe17;
input 	dffe162;
output 	dffe163;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[15]~q ;
wire \xordvalue[10]~q ;
wire \Add0~1_sumout ;
wire \a[14]~q ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \a[13]~q ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \a[12]~q ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \a[11]~q ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \a[10]~q ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \a[9]~q ;
wire \xordvalue[0]~q ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \a[8]~q ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \a[7]~q ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \a[6]~q ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \a[5]~q ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \a[4]~q ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \a[3]~q ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~51 ;
wire \a[2]~q ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~55 ;
wire \a[1]~q ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~59 ;
wire \a[0]~q ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~63 ;


nco_test_lpm_add_sub_38 u0(
	.a_15(\a[15]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.a_14(\a[14]~q ),
	.a_13(\a[13]~q ),
	.a_12(\a[12]~q ),
	.a_11(\a[11]~q ),
	.a_10(\a[10]~q ),
	.a_9(\a[9]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_8(\a[8]~q ),
	.a_7(\a[7]~q ),
	.a_6(\a[6]~q ),
	.a_5(\a[5]~q ),
	.a_4(\a[4]~q ),
	.a_3(\a[3]~q ),
	.a_2(\a[2]~q ),
	.a_1(\a[1]~q ),
	.a_0(\a[0]~q ),
	.dffe16(dffe16),
	.dffe15(dffe15),
	.dffe14(dffe14),
	.dffe13(dffe13),
	.dffe12(dffe12),
	.dffe11(dffe11),
	.dffe10(dffe10),
	.dffe9(dffe9),
	.dffe8(dffe8),
	.dffe7(dffe7),
	.dffe6(dffe6),
	.dffe5(dffe5),
	.dffe4(dffe4),
	.dffe3(dffe3),
	.dffe2(dffe2),
	.dffe1(dffe1),
	.dffe161(dffe163),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(dffe161),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "on";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~5 .shared_arith = "on";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~9 .shared_arith = "on";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~13 .shared_arith = "on";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~17 .shared_arith = "on";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "on";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(dffe162),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~25 .shared_arith = "on";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~29 .shared_arith = "on";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~33 .shared_arith = "on";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~37 .shared_arith = "on";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(\Add0~47 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~41 .shared_arith = "on";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(\Add0~51 ),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout(\Add0~47 ));
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~45 .shared_arith = "on";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(\Add0~55 ),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout(\Add0~51 ));
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~49 .shared_arith = "on";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(\Add0~59 ),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout(\Add0~55 ));
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~53 .shared_arith = "on";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(\Add0~63 ),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout(\Add0~59 ));
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~57 .shared_arith = "on";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!dffe17),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout(\Add0~63 ));
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add0~61 .shared_arith = "on";

endmodule

module nco_test_lpm_add_sub_38 (
	a_15,
	xordvalue_10,
	a_14,
	a_13,
	a_12,
	a_11,
	a_10,
	a_9,
	xordvalue_0,
	a_8,
	a_7,
	a_6,
	a_5,
	a_4,
	a_3,
	a_2,
	a_1,
	a_0,
	dffe16,
	dffe15,
	dffe14,
	dffe13,
	dffe12,
	dffe11,
	dffe10,
	dffe9,
	dffe8,
	dffe7,
	dffe6,
	dffe5,
	dffe4,
	dffe3,
	dffe2,
	dffe1,
	dffe161,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_15;
input 	xordvalue_10;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_10;
input 	a_9;
input 	xordvalue_0;
input 	a_8;
input 	a_7;
input 	a_6;
input 	a_5;
input 	a_4;
input 	a_3;
input 	a_2;
input 	a_1;
input 	a_0;
output 	dffe16;
output 	dffe15;
output 	dffe14;
output 	dffe13;
output 	dffe12;
output 	dffe11;
output 	dffe10;
output 	dffe9;
output 	dffe8;
output 	dffe7;
output 	dffe6;
output 	dffe5;
output 	dffe4;
output 	dffe3;
output 	dffe2;
output 	dffe1;
output 	dffe161;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_add_sub_hdg_2 auto_generated(
	.a_15(a_15),
	.xordvalue_10(xordvalue_10),
	.a_14(a_14),
	.a_13(a_13),
	.a_12(a_12),
	.a_11(a_11),
	.a_10(a_10),
	.a_9(a_9),
	.xordvalue_0(xordvalue_0),
	.a_8(a_8),
	.a_7(a_7),
	.a_6(a_6),
	.a_5(a_5),
	.a_4(a_4),
	.a_3(a_3),
	.a_2(a_2),
	.a_1(a_1),
	.a_0(a_0),
	.dffe161(dffe16),
	.dffe151(dffe15),
	.dffe141(dffe14),
	.dffe131(dffe13),
	.dffe121(dffe12),
	.dffe111(dffe11),
	.dffe101(dffe10),
	.dffe91(dffe9),
	.dffe81(dffe8),
	.dffe71(dffe7),
	.dffe61(dffe6),
	.dffe51(dffe5),
	.dffe41(dffe4),
	.dffe31(dffe3),
	.dffe21(dffe2),
	.dffe17(dffe1),
	.dffe162(dffe161),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module nco_test_add_sub_hdg_2 (
	a_15,
	xordvalue_10,
	a_14,
	a_13,
	a_12,
	a_11,
	a_10,
	a_9,
	xordvalue_0,
	a_8,
	a_7,
	a_6,
	a_5,
	a_4,
	a_3,
	a_2,
	a_1,
	a_0,
	dffe161,
	dffe151,
	dffe141,
	dffe131,
	dffe121,
	dffe111,
	dffe101,
	dffe91,
	dffe81,
	dffe71,
	dffe61,
	dffe51,
	dffe41,
	dffe31,
	dffe21,
	dffe17,
	dffe162,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_15;
input 	xordvalue_10;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_10;
input 	a_9;
input 	xordvalue_0;
input 	a_8;
input 	a_7;
input 	a_6;
input 	a_5;
input 	a_4;
input 	a_3;
input 	a_2;
input 	a_1;
input 	a_0;
output 	dffe161;
output 	dffe151;
output 	dffe141;
output 	dffe131;
output 	dffe121;
output 	dffe111;
output 	dffe101;
output 	dffe91;
output 	dffe81;
output 	dffe71;
output 	dffe61;
output 	dffe51;
output 	dffe41;
output 	dffe31;
output 	dffe21;
output 	dffe17;
output 	dffe162;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~COUT ;
wire \add_sub_cella[12]~COUT ;
wire \add_sub_cella[13]~COUT ;
wire \add_sub_cella[14]~COUT ;
wire \add_sub_cella[15]~sumout ;
wire \add_sub_cella[14]~sumout ;
wire \add_sub_cella[13]~sumout ;
wire \add_sub_cella[12]~sumout ;
wire \add_sub_cella[11]~sumout ;
wire \add_sub_cella[10]~sumout ;
wire \add_sub_cella[9]~sumout ;
wire \add_sub_cella[8]~sumout ;
wire \add_sub_cella[7]~sumout ;
wire \add_sub_cella[6]~sumout ;
wire \add_sub_cella[5]~sumout ;
wire \add_sub_cella[4]~sumout ;
wire \add_sub_cella[3]~sumout ;
wire \add_sub_cella[2]~sumout ;
wire \add_sub_cella[1]~sumout ;
wire \add_sub_cella[0]~sumout ;


dffeas dffe16(
	.clk(clock),
	.d(\add_sub_cella[15]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe161),
	.prn(vcc));
defparam dffe16.is_wysiwyg = "true";
defparam dffe16.power_up = "low";

dffeas dffe15(
	.clk(clock),
	.d(\add_sub_cella[14]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe151),
	.prn(vcc));
defparam dffe15.is_wysiwyg = "true";
defparam dffe15.power_up = "low";

dffeas dffe14(
	.clk(clock),
	.d(\add_sub_cella[13]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe141),
	.prn(vcc));
defparam dffe14.is_wysiwyg = "true";
defparam dffe14.power_up = "low";

dffeas dffe13(
	.clk(clock),
	.d(\add_sub_cella[12]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe131),
	.prn(vcc));
defparam dffe13.is_wysiwyg = "true";
defparam dffe13.power_up = "low";

dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe17),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

arriav_lcell_comb \dffe16~_wirecell (
	.dataa(!dffe161),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(dffe162),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffe16~_wirecell .extended_lut = "off";
defparam \dffe16~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dffe16~_wirecell .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(\add_sub_cella[11]~COUT ),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[12] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[11]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[12]~sumout ),
	.cout(\add_sub_cella[12]~COUT ),
	.shareout());
defparam \add_sub_cella[12] .extended_lut = "off";
defparam \add_sub_cella[12] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[12] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[13] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[12]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[13]~sumout ),
	.cout(\add_sub_cella[13]~COUT ),
	.shareout());
defparam \add_sub_cella[13] .extended_lut = "off";
defparam \add_sub_cella[13] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[13] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[14] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[13]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[14]~sumout ),
	.cout(\add_sub_cella[14]~COUT ),
	.shareout());
defparam \add_sub_cella[14] .extended_lut = "off";
defparam \add_sub_cella[14] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[14] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[15] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[14]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[15]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[15] .extended_lut = "off";
defparam \add_sub_cella[15] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[15] .shared_arith = "off";

endmodule

module nco_test_cordic_zxor_1p_lpm_3 (
	sin_o_0,
	dffe16,
	dffe15,
	dffe14,
	dffe161,
	dffe13,
	dffe12,
	dffe151,
	dffe11,
	dffe141,
	dffe10,
	dffe131,
	dffe9,
	dffe121,
	dffe8,
	dffe111,
	dffe7,
	dffe101,
	dffe6,
	dffe91,
	dffe5,
	dffe81,
	dffe4,
	dffe71,
	dffe3,
	dffe61,
	dffe2,
	dffe51,
	dffe1,
	dffe41,
	dffe31,
	dffe21,
	dffe17,
	dffe162,
	dffe163,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	sin_o_0;
output 	dffe16;
output 	dffe15;
output 	dffe14;
input 	dffe161;
output 	dffe13;
output 	dffe12;
input 	dffe151;
output 	dffe11;
input 	dffe141;
output 	dffe10;
input 	dffe131;
output 	dffe9;
input 	dffe121;
output 	dffe8;
input 	dffe111;
output 	dffe7;
input 	dffe101;
output 	dffe6;
input 	dffe91;
output 	dffe5;
input 	dffe81;
output 	dffe4;
input 	dffe71;
output 	dffe3;
input 	dffe61;
output 	dffe2;
input 	dffe51;
output 	dffe1;
input 	dffe41;
input 	dffe31;
input 	dffe21;
input 	dffe17;
input 	dffe162;
output 	dffe163;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[15]~q ;
wire \xordvalue[10]~q ;
wire \Add0~1_sumout ;
wire \a[14]~q ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \a[13]~q ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \a[12]~q ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \a[11]~q ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \a[10]~q ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \a[9]~q ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \a[8]~q ;
wire \xordvalue[0]~q ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \a[7]~q ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \a[6]~q ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \a[5]~q ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \a[4]~q ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \a[3]~q ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~51 ;
wire \a[2]~q ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~55 ;
wire \a[1]~q ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~59 ;
wire \a[0]~q ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~63 ;


nco_test_lpm_add_sub_39 u0(
	.a_15(\a[15]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.a_14(\a[14]~q ),
	.a_13(\a[13]~q ),
	.a_12(\a[12]~q ),
	.a_11(\a[11]~q ),
	.a_10(\a[10]~q ),
	.a_9(\a[9]~q ),
	.a_8(\a[8]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_7(\a[7]~q ),
	.a_6(\a[6]~q ),
	.a_5(\a[5]~q ),
	.a_4(\a[4]~q ),
	.a_3(\a[3]~q ),
	.a_2(\a[2]~q ),
	.a_1(\a[1]~q ),
	.a_0(\a[0]~q ),
	.dffe16(dffe16),
	.dffe15(dffe15),
	.dffe14(dffe14),
	.dffe13(dffe13),
	.dffe12(dffe12),
	.dffe11(dffe11),
	.dffe10(dffe10),
	.dffe9(dffe9),
	.dffe8(dffe8),
	.dffe7(dffe7),
	.dffe6(dffe6),
	.dffe5(dffe5),
	.dffe4(dffe4),
	.dffe3(dffe3),
	.dffe2(dffe2),
	.dffe1(dffe1),
	.dffe161(dffe163),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(dffe161),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "on";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~5 .shared_arith = "on";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~9 .shared_arith = "on";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~13 .shared_arith = "on";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~17 .shared_arith = "on";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "on";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~25 .shared_arith = "on";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(dffe162),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~29 .shared_arith = "on";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~33 .shared_arith = "on";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~37 .shared_arith = "on";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(\Add0~47 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~41 .shared_arith = "on";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(\Add0~51 ),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout(\Add0~47 ));
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~45 .shared_arith = "on";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(\Add0~55 ),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout(\Add0~51 ));
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~49 .shared_arith = "on";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(\Add0~59 ),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout(\Add0~55 ));
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~53 .shared_arith = "on";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(\Add0~63 ),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout(\Add0~59 ));
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~57 .shared_arith = "on";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!dffe17),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout(\Add0~63 ));
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add0~61 .shared_arith = "on";

endmodule

module nco_test_lpm_add_sub_39 (
	a_15,
	xordvalue_10,
	a_14,
	a_13,
	a_12,
	a_11,
	a_10,
	a_9,
	a_8,
	xordvalue_0,
	a_7,
	a_6,
	a_5,
	a_4,
	a_3,
	a_2,
	a_1,
	a_0,
	dffe16,
	dffe15,
	dffe14,
	dffe13,
	dffe12,
	dffe11,
	dffe10,
	dffe9,
	dffe8,
	dffe7,
	dffe6,
	dffe5,
	dffe4,
	dffe3,
	dffe2,
	dffe1,
	dffe161,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_15;
input 	xordvalue_10;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_10;
input 	a_9;
input 	a_8;
input 	xordvalue_0;
input 	a_7;
input 	a_6;
input 	a_5;
input 	a_4;
input 	a_3;
input 	a_2;
input 	a_1;
input 	a_0;
output 	dffe16;
output 	dffe15;
output 	dffe14;
output 	dffe13;
output 	dffe12;
output 	dffe11;
output 	dffe10;
output 	dffe9;
output 	dffe8;
output 	dffe7;
output 	dffe6;
output 	dffe5;
output 	dffe4;
output 	dffe3;
output 	dffe2;
output 	dffe1;
output 	dffe161;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_add_sub_hdg_3 auto_generated(
	.a_15(a_15),
	.xordvalue_10(xordvalue_10),
	.a_14(a_14),
	.a_13(a_13),
	.a_12(a_12),
	.a_11(a_11),
	.a_10(a_10),
	.a_9(a_9),
	.a_8(a_8),
	.xordvalue_0(xordvalue_0),
	.a_7(a_7),
	.a_6(a_6),
	.a_5(a_5),
	.a_4(a_4),
	.a_3(a_3),
	.a_2(a_2),
	.a_1(a_1),
	.a_0(a_0),
	.dffe161(dffe16),
	.dffe151(dffe15),
	.dffe141(dffe14),
	.dffe131(dffe13),
	.dffe121(dffe12),
	.dffe111(dffe11),
	.dffe101(dffe10),
	.dffe91(dffe9),
	.dffe81(dffe8),
	.dffe71(dffe7),
	.dffe61(dffe6),
	.dffe51(dffe5),
	.dffe41(dffe4),
	.dffe31(dffe3),
	.dffe21(dffe2),
	.dffe17(dffe1),
	.dffe162(dffe161),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module nco_test_add_sub_hdg_3 (
	a_15,
	xordvalue_10,
	a_14,
	a_13,
	a_12,
	a_11,
	a_10,
	a_9,
	a_8,
	xordvalue_0,
	a_7,
	a_6,
	a_5,
	a_4,
	a_3,
	a_2,
	a_1,
	a_0,
	dffe161,
	dffe151,
	dffe141,
	dffe131,
	dffe121,
	dffe111,
	dffe101,
	dffe91,
	dffe81,
	dffe71,
	dffe61,
	dffe51,
	dffe41,
	dffe31,
	dffe21,
	dffe17,
	dffe162,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_15;
input 	xordvalue_10;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_10;
input 	a_9;
input 	a_8;
input 	xordvalue_0;
input 	a_7;
input 	a_6;
input 	a_5;
input 	a_4;
input 	a_3;
input 	a_2;
input 	a_1;
input 	a_0;
output 	dffe161;
output 	dffe151;
output 	dffe141;
output 	dffe131;
output 	dffe121;
output 	dffe111;
output 	dffe101;
output 	dffe91;
output 	dffe81;
output 	dffe71;
output 	dffe61;
output 	dffe51;
output 	dffe41;
output 	dffe31;
output 	dffe21;
output 	dffe17;
output 	dffe162;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~COUT ;
wire \add_sub_cella[12]~COUT ;
wire \add_sub_cella[13]~COUT ;
wire \add_sub_cella[14]~COUT ;
wire \add_sub_cella[15]~sumout ;
wire \add_sub_cella[14]~sumout ;
wire \add_sub_cella[13]~sumout ;
wire \add_sub_cella[12]~sumout ;
wire \add_sub_cella[11]~sumout ;
wire \add_sub_cella[10]~sumout ;
wire \add_sub_cella[9]~sumout ;
wire \add_sub_cella[8]~sumout ;
wire \add_sub_cella[7]~sumout ;
wire \add_sub_cella[6]~sumout ;
wire \add_sub_cella[5]~sumout ;
wire \add_sub_cella[4]~sumout ;
wire \add_sub_cella[3]~sumout ;
wire \add_sub_cella[2]~sumout ;
wire \add_sub_cella[1]~sumout ;
wire \add_sub_cella[0]~sumout ;


dffeas dffe16(
	.clk(clock),
	.d(\add_sub_cella[15]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe161),
	.prn(vcc));
defparam dffe16.is_wysiwyg = "true";
defparam dffe16.power_up = "low";

dffeas dffe15(
	.clk(clock),
	.d(\add_sub_cella[14]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe151),
	.prn(vcc));
defparam dffe15.is_wysiwyg = "true";
defparam dffe15.power_up = "low";

dffeas dffe14(
	.clk(clock),
	.d(\add_sub_cella[13]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe141),
	.prn(vcc));
defparam dffe14.is_wysiwyg = "true";
defparam dffe14.power_up = "low";

dffeas dffe13(
	.clk(clock),
	.d(\add_sub_cella[12]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe131),
	.prn(vcc));
defparam dffe13.is_wysiwyg = "true";
defparam dffe13.power_up = "low";

dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe17),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

arriav_lcell_comb \dffe16~_wirecell (
	.dataa(!dffe161),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(dffe162),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffe16~_wirecell .extended_lut = "off";
defparam \dffe16~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dffe16~_wirecell .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(\add_sub_cella[11]~COUT ),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[12] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[11]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[12]~sumout ),
	.cout(\add_sub_cella[12]~COUT ),
	.shareout());
defparam \add_sub_cella[12] .extended_lut = "off";
defparam \add_sub_cella[12] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[12] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[13] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[12]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[13]~sumout ),
	.cout(\add_sub_cella[13]~COUT ),
	.shareout());
defparam \add_sub_cella[13] .extended_lut = "off";
defparam \add_sub_cella[13] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[13] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[14] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[13]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[14]~sumout ),
	.cout(\add_sub_cella[14]~COUT ),
	.shareout());
defparam \add_sub_cella[14] .extended_lut = "off";
defparam \add_sub_cella[14] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[14] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[15] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[14]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[15]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[15] .extended_lut = "off";
defparam \add_sub_cella[15] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[15] .shared_arith = "off";

endmodule

module nco_test_cordic_zxor_1p_lpm_4 (
	sin_o_0,
	dffe16,
	dffe15,
	dffe14,
	dffe161,
	dffe13,
	dffe12,
	dffe151,
	dffe11,
	dffe141,
	dffe10,
	dffe131,
	dffe9,
	dffe121,
	dffe8,
	dffe111,
	dffe7,
	dffe101,
	dffe6,
	dffe91,
	dffe5,
	dffe81,
	dffe4,
	dffe71,
	dffe3,
	dffe61,
	dffe2,
	dffe51,
	dffe1,
	dffe41,
	dffe31,
	dffe21,
	dffe17,
	dffe162,
	dffe163,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	sin_o_0;
output 	dffe16;
output 	dffe15;
output 	dffe14;
input 	dffe161;
output 	dffe13;
output 	dffe12;
input 	dffe151;
output 	dffe11;
input 	dffe141;
output 	dffe10;
input 	dffe131;
output 	dffe9;
input 	dffe121;
output 	dffe8;
input 	dffe111;
output 	dffe7;
input 	dffe101;
output 	dffe6;
input 	dffe91;
output 	dffe5;
input 	dffe81;
output 	dffe4;
input 	dffe71;
output 	dffe3;
input 	dffe61;
output 	dffe2;
input 	dffe51;
output 	dffe1;
input 	dffe41;
input 	dffe31;
input 	dffe21;
input 	dffe17;
input 	dffe162;
output 	dffe163;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[15]~q ;
wire \xordvalue[0]~q ;
wire \Add0~1_sumout ;
wire \a[14]~q ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \a[13]~q ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \a[12]~q ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \a[11]~q ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \a[10]~q ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \a[9]~q ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \a[8]~q ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \a[7]~q ;
wire \xordvalue[1]~q ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \a[6]~q ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \a[5]~q ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \a[4]~q ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \a[3]~q ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~51 ;
wire \a[2]~q ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~55 ;
wire \a[1]~q ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~59 ;
wire \a[0]~q ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~63 ;


nco_test_lpm_add_sub_40 u0(
	.a_15(\a[15]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_14(\a[14]~q ),
	.a_13(\a[13]~q ),
	.a_12(\a[12]~q ),
	.a_11(\a[11]~q ),
	.a_10(\a[10]~q ),
	.a_9(\a[9]~q ),
	.a_8(\a[8]~q ),
	.a_7(\a[7]~q ),
	.xordvalue_1(\xordvalue[1]~q ),
	.a_6(\a[6]~q ),
	.a_5(\a[5]~q ),
	.a_4(\a[4]~q ),
	.a_3(\a[3]~q ),
	.a_2(\a[2]~q ),
	.a_1(\a[1]~q ),
	.a_0(\a[0]~q ),
	.dffe16(dffe16),
	.dffe15(dffe15),
	.dffe14(dffe14),
	.dffe13(dffe13),
	.dffe12(dffe12),
	.dffe11(dffe11),
	.dffe10(dffe10),
	.dffe9(dffe9),
	.dffe8(dffe8),
	.dffe7(dffe7),
	.dffe6(dffe6),
	.dffe5(dffe5),
	.dffe4(dffe4),
	.dffe3(dffe3),
	.dffe2(dffe2),
	.dffe1(dffe1),
	.dffe161(dffe163),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(dffe161),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "on";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~5 .shared_arith = "on";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~9 .shared_arith = "on";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~13 .shared_arith = "on";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~17 .shared_arith = "on";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "on";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~25 .shared_arith = "on";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~29 .shared_arith = "on";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \xordvalue[1] (
	.clk(clk),
	.d(dffe162),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[1]~q ),
	.prn(vcc));
defparam \xordvalue[1] .is_wysiwyg = "true";
defparam \xordvalue[1] .power_up = "low";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~33 .shared_arith = "on";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~37 .shared_arith = "on";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(\Add0~47 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~41 .shared_arith = "on";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(\Add0~51 ),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout(\Add0~47 ));
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~45 .shared_arith = "on";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(\Add0~55 ),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout(\Add0~51 ));
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~49 .shared_arith = "on";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(\Add0~59 ),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout(\Add0~55 ));
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~53 .shared_arith = "on";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(\Add0~63 ),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout(\Add0~59 ));
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~57 .shared_arith = "on";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!dffe17),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout(\Add0~63 ));
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add0~61 .shared_arith = "on";

endmodule

module nco_test_lpm_add_sub_40 (
	a_15,
	xordvalue_0,
	a_14,
	a_13,
	a_12,
	a_11,
	a_10,
	a_9,
	a_8,
	a_7,
	xordvalue_1,
	a_6,
	a_5,
	a_4,
	a_3,
	a_2,
	a_1,
	a_0,
	dffe16,
	dffe15,
	dffe14,
	dffe13,
	dffe12,
	dffe11,
	dffe10,
	dffe9,
	dffe8,
	dffe7,
	dffe6,
	dffe5,
	dffe4,
	dffe3,
	dffe2,
	dffe1,
	dffe161,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_15;
input 	xordvalue_0;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_10;
input 	a_9;
input 	a_8;
input 	a_7;
input 	xordvalue_1;
input 	a_6;
input 	a_5;
input 	a_4;
input 	a_3;
input 	a_2;
input 	a_1;
input 	a_0;
output 	dffe16;
output 	dffe15;
output 	dffe14;
output 	dffe13;
output 	dffe12;
output 	dffe11;
output 	dffe10;
output 	dffe9;
output 	dffe8;
output 	dffe7;
output 	dffe6;
output 	dffe5;
output 	dffe4;
output 	dffe3;
output 	dffe2;
output 	dffe1;
output 	dffe161;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_add_sub_hdg_4 auto_generated(
	.a_15(a_15),
	.xordvalue_0(xordvalue_0),
	.a_14(a_14),
	.a_13(a_13),
	.a_12(a_12),
	.a_11(a_11),
	.a_10(a_10),
	.a_9(a_9),
	.a_8(a_8),
	.a_7(a_7),
	.xordvalue_1(xordvalue_1),
	.a_6(a_6),
	.a_5(a_5),
	.a_4(a_4),
	.a_3(a_3),
	.a_2(a_2),
	.a_1(a_1),
	.a_0(a_0),
	.dffe161(dffe16),
	.dffe151(dffe15),
	.dffe141(dffe14),
	.dffe131(dffe13),
	.dffe121(dffe12),
	.dffe111(dffe11),
	.dffe101(dffe10),
	.dffe91(dffe9),
	.dffe81(dffe8),
	.dffe71(dffe7),
	.dffe61(dffe6),
	.dffe51(dffe5),
	.dffe41(dffe4),
	.dffe31(dffe3),
	.dffe21(dffe2),
	.dffe17(dffe1),
	.dffe162(dffe161),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module nco_test_add_sub_hdg_4 (
	a_15,
	xordvalue_0,
	a_14,
	a_13,
	a_12,
	a_11,
	a_10,
	a_9,
	a_8,
	a_7,
	xordvalue_1,
	a_6,
	a_5,
	a_4,
	a_3,
	a_2,
	a_1,
	a_0,
	dffe161,
	dffe151,
	dffe141,
	dffe131,
	dffe121,
	dffe111,
	dffe101,
	dffe91,
	dffe81,
	dffe71,
	dffe61,
	dffe51,
	dffe41,
	dffe31,
	dffe21,
	dffe17,
	dffe162,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_15;
input 	xordvalue_0;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_10;
input 	a_9;
input 	a_8;
input 	a_7;
input 	xordvalue_1;
input 	a_6;
input 	a_5;
input 	a_4;
input 	a_3;
input 	a_2;
input 	a_1;
input 	a_0;
output 	dffe161;
output 	dffe151;
output 	dffe141;
output 	dffe131;
output 	dffe121;
output 	dffe111;
output 	dffe101;
output 	dffe91;
output 	dffe81;
output 	dffe71;
output 	dffe61;
output 	dffe51;
output 	dffe41;
output 	dffe31;
output 	dffe21;
output 	dffe17;
output 	dffe162;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~COUT ;
wire \add_sub_cella[12]~COUT ;
wire \add_sub_cella[13]~COUT ;
wire \add_sub_cella[14]~COUT ;
wire \add_sub_cella[15]~sumout ;
wire \add_sub_cella[14]~sumout ;
wire \add_sub_cella[13]~sumout ;
wire \add_sub_cella[12]~sumout ;
wire \add_sub_cella[11]~sumout ;
wire \add_sub_cella[10]~sumout ;
wire \add_sub_cella[9]~sumout ;
wire \add_sub_cella[8]~sumout ;
wire \add_sub_cella[7]~sumout ;
wire \add_sub_cella[6]~sumout ;
wire \add_sub_cella[5]~sumout ;
wire \add_sub_cella[4]~sumout ;
wire \add_sub_cella[3]~sumout ;
wire \add_sub_cella[2]~sumout ;
wire \add_sub_cella[1]~sumout ;
wire \add_sub_cella[0]~sumout ;


dffeas dffe16(
	.clk(clock),
	.d(\add_sub_cella[15]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe161),
	.prn(vcc));
defparam dffe16.is_wysiwyg = "true";
defparam dffe16.power_up = "low";

dffeas dffe15(
	.clk(clock),
	.d(\add_sub_cella[14]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe151),
	.prn(vcc));
defparam dffe15.is_wysiwyg = "true";
defparam dffe15.power_up = "low";

dffeas dffe14(
	.clk(clock),
	.d(\add_sub_cella[13]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe141),
	.prn(vcc));
defparam dffe14.is_wysiwyg = "true";
defparam dffe14.power_up = "low";

dffeas dffe13(
	.clk(clock),
	.d(\add_sub_cella[12]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe131),
	.prn(vcc));
defparam dffe13.is_wysiwyg = "true";
defparam dffe13.power_up = "low";

dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe17),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

arriav_lcell_comb \dffe16~_wirecell (
	.dataa(!dffe161),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(dffe162),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffe16~_wirecell .extended_lut = "off";
defparam \dffe16~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dffe16~_wirecell .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_1),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_1),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_1),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(\add_sub_cella[11]~COUT ),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[12] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[11]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[12]~sumout ),
	.cout(\add_sub_cella[12]~COUT ),
	.shareout());
defparam \add_sub_cella[12] .extended_lut = "off";
defparam \add_sub_cella[12] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[12] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[13] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[12]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[13]~sumout ),
	.cout(\add_sub_cella[13]~COUT ),
	.shareout());
defparam \add_sub_cella[13] .extended_lut = "off";
defparam \add_sub_cella[13] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[13] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[14] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[13]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[14]~sumout ),
	.cout(\add_sub_cella[14]~COUT ),
	.shareout());
defparam \add_sub_cella[14] .extended_lut = "off";
defparam \add_sub_cella[14] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[14] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[15] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[14]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[15]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[15] .extended_lut = "off";
defparam \add_sub_cella[15] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[15] .shared_arith = "off";

endmodule

module nco_test_cordic_zxor_1p_lpm_5 (
	sin_o_0,
	dffe16,
	dffe15,
	dffe14,
	dffe161,
	dffe13,
	dffe12,
	dffe151,
	dffe11,
	dffe141,
	dffe10,
	dffe131,
	dffe9,
	dffe121,
	dffe8,
	dffe111,
	dffe7,
	dffe101,
	dffe6,
	dffe91,
	dffe5,
	dffe81,
	dffe4,
	dffe71,
	dffe3,
	dffe61,
	dffe2,
	dffe51,
	dffe1,
	dffe41,
	dffe31,
	dffe21,
	dffe17,
	dffe162,
	dffe163,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	sin_o_0;
output 	dffe16;
output 	dffe15;
output 	dffe14;
input 	dffe161;
output 	dffe13;
output 	dffe12;
input 	dffe151;
output 	dffe11;
input 	dffe141;
output 	dffe10;
input 	dffe131;
output 	dffe9;
input 	dffe121;
output 	dffe8;
input 	dffe111;
output 	dffe7;
input 	dffe101;
output 	dffe6;
input 	dffe91;
output 	dffe5;
input 	dffe81;
output 	dffe4;
input 	dffe71;
output 	dffe3;
input 	dffe61;
output 	dffe2;
input 	dffe51;
output 	dffe1;
input 	dffe41;
input 	dffe31;
input 	dffe21;
input 	dffe17;
input 	dffe162;
output 	dffe163;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[15]~q ;
wire \xordvalue[10]~q ;
wire \Add0~1_sumout ;
wire \a[14]~q ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \a[13]~q ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \a[12]~q ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \a[11]~q ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \a[10]~q ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \a[9]~q ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \a[8]~q ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \a[7]~q ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \a[6]~q ;
wire \xordvalue[0]~q ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \a[5]~q ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \a[4]~q ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \a[3]~q ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~51 ;
wire \a[2]~q ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~55 ;
wire \a[1]~q ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~59 ;
wire \a[0]~q ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~63 ;


nco_test_lpm_add_sub_41 u0(
	.a_15(\a[15]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.a_14(\a[14]~q ),
	.a_13(\a[13]~q ),
	.a_12(\a[12]~q ),
	.a_11(\a[11]~q ),
	.a_10(\a[10]~q ),
	.a_9(\a[9]~q ),
	.a_8(\a[8]~q ),
	.a_7(\a[7]~q ),
	.a_6(\a[6]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_5(\a[5]~q ),
	.a_4(\a[4]~q ),
	.a_3(\a[3]~q ),
	.a_2(\a[2]~q ),
	.a_1(\a[1]~q ),
	.a_0(\a[0]~q ),
	.dffe16(dffe16),
	.dffe15(dffe15),
	.dffe14(dffe14),
	.dffe13(dffe13),
	.dffe12(dffe12),
	.dffe11(dffe11),
	.dffe10(dffe10),
	.dffe9(dffe9),
	.dffe8(dffe8),
	.dffe7(dffe7),
	.dffe6(dffe6),
	.dffe5(dffe5),
	.dffe4(dffe4),
	.dffe3(dffe3),
	.dffe2(dffe2),
	.dffe1(dffe1),
	.dffe161(dffe163),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(dffe161),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "on";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~5 .shared_arith = "on";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~9 .shared_arith = "on";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~13 .shared_arith = "on";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~17 .shared_arith = "on";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "on";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~25 .shared_arith = "on";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~29 .shared_arith = "on";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~33 .shared_arith = "on";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(dffe162),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~37 .shared_arith = "on";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(\Add0~47 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~41 .shared_arith = "on";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(\Add0~51 ),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout(\Add0~47 ));
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~45 .shared_arith = "on";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(\Add0~55 ),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout(\Add0~51 ));
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~49 .shared_arith = "on";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(\Add0~59 ),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout(\Add0~55 ));
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~53 .shared_arith = "on";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(\Add0~63 ),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout(\Add0~59 ));
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~57 .shared_arith = "on";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!dffe17),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout(\Add0~63 ));
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add0~61 .shared_arith = "on";

endmodule

module nco_test_lpm_add_sub_41 (
	a_15,
	xordvalue_10,
	a_14,
	a_13,
	a_12,
	a_11,
	a_10,
	a_9,
	a_8,
	a_7,
	a_6,
	xordvalue_0,
	a_5,
	a_4,
	a_3,
	a_2,
	a_1,
	a_0,
	dffe16,
	dffe15,
	dffe14,
	dffe13,
	dffe12,
	dffe11,
	dffe10,
	dffe9,
	dffe8,
	dffe7,
	dffe6,
	dffe5,
	dffe4,
	dffe3,
	dffe2,
	dffe1,
	dffe161,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_15;
input 	xordvalue_10;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_10;
input 	a_9;
input 	a_8;
input 	a_7;
input 	a_6;
input 	xordvalue_0;
input 	a_5;
input 	a_4;
input 	a_3;
input 	a_2;
input 	a_1;
input 	a_0;
output 	dffe16;
output 	dffe15;
output 	dffe14;
output 	dffe13;
output 	dffe12;
output 	dffe11;
output 	dffe10;
output 	dffe9;
output 	dffe8;
output 	dffe7;
output 	dffe6;
output 	dffe5;
output 	dffe4;
output 	dffe3;
output 	dffe2;
output 	dffe1;
output 	dffe161;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_add_sub_hdg_5 auto_generated(
	.a_15(a_15),
	.xordvalue_10(xordvalue_10),
	.a_14(a_14),
	.a_13(a_13),
	.a_12(a_12),
	.a_11(a_11),
	.a_10(a_10),
	.a_9(a_9),
	.a_8(a_8),
	.a_7(a_7),
	.a_6(a_6),
	.xordvalue_0(xordvalue_0),
	.a_5(a_5),
	.a_4(a_4),
	.a_3(a_3),
	.a_2(a_2),
	.a_1(a_1),
	.a_0(a_0),
	.dffe161(dffe16),
	.dffe151(dffe15),
	.dffe141(dffe14),
	.dffe131(dffe13),
	.dffe121(dffe12),
	.dffe111(dffe11),
	.dffe101(dffe10),
	.dffe91(dffe9),
	.dffe81(dffe8),
	.dffe71(dffe7),
	.dffe61(dffe6),
	.dffe51(dffe5),
	.dffe41(dffe4),
	.dffe31(dffe3),
	.dffe21(dffe2),
	.dffe17(dffe1),
	.dffe162(dffe161),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module nco_test_add_sub_hdg_5 (
	a_15,
	xordvalue_10,
	a_14,
	a_13,
	a_12,
	a_11,
	a_10,
	a_9,
	a_8,
	a_7,
	a_6,
	xordvalue_0,
	a_5,
	a_4,
	a_3,
	a_2,
	a_1,
	a_0,
	dffe161,
	dffe151,
	dffe141,
	dffe131,
	dffe121,
	dffe111,
	dffe101,
	dffe91,
	dffe81,
	dffe71,
	dffe61,
	dffe51,
	dffe41,
	dffe31,
	dffe21,
	dffe17,
	dffe162,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_15;
input 	xordvalue_10;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_10;
input 	a_9;
input 	a_8;
input 	a_7;
input 	a_6;
input 	xordvalue_0;
input 	a_5;
input 	a_4;
input 	a_3;
input 	a_2;
input 	a_1;
input 	a_0;
output 	dffe161;
output 	dffe151;
output 	dffe141;
output 	dffe131;
output 	dffe121;
output 	dffe111;
output 	dffe101;
output 	dffe91;
output 	dffe81;
output 	dffe71;
output 	dffe61;
output 	dffe51;
output 	dffe41;
output 	dffe31;
output 	dffe21;
output 	dffe17;
output 	dffe162;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~COUT ;
wire \add_sub_cella[12]~COUT ;
wire \add_sub_cella[13]~COUT ;
wire \add_sub_cella[14]~COUT ;
wire \add_sub_cella[15]~sumout ;
wire \add_sub_cella[14]~sumout ;
wire \add_sub_cella[13]~sumout ;
wire \add_sub_cella[12]~sumout ;
wire \add_sub_cella[11]~sumout ;
wire \add_sub_cella[10]~sumout ;
wire \add_sub_cella[9]~sumout ;
wire \add_sub_cella[8]~sumout ;
wire \add_sub_cella[7]~sumout ;
wire \add_sub_cella[6]~sumout ;
wire \add_sub_cella[5]~sumout ;
wire \add_sub_cella[4]~sumout ;
wire \add_sub_cella[3]~sumout ;
wire \add_sub_cella[2]~sumout ;
wire \add_sub_cella[1]~sumout ;
wire \add_sub_cella[0]~sumout ;


dffeas dffe16(
	.clk(clock),
	.d(\add_sub_cella[15]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe161),
	.prn(vcc));
defparam dffe16.is_wysiwyg = "true";
defparam dffe16.power_up = "low";

dffeas dffe15(
	.clk(clock),
	.d(\add_sub_cella[14]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe151),
	.prn(vcc));
defparam dffe15.is_wysiwyg = "true";
defparam dffe15.power_up = "low";

dffeas dffe14(
	.clk(clock),
	.d(\add_sub_cella[13]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe141),
	.prn(vcc));
defparam dffe14.is_wysiwyg = "true";
defparam dffe14.power_up = "low";

dffeas dffe13(
	.clk(clock),
	.d(\add_sub_cella[12]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe131),
	.prn(vcc));
defparam dffe13.is_wysiwyg = "true";
defparam dffe13.power_up = "low";

dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe17),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

arriav_lcell_comb \dffe16~_wirecell (
	.dataa(!dffe161),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(dffe162),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffe16~_wirecell .extended_lut = "off";
defparam \dffe16~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dffe16~_wirecell .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(\add_sub_cella[11]~COUT ),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[12] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[11]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[12]~sumout ),
	.cout(\add_sub_cella[12]~COUT ),
	.shareout());
defparam \add_sub_cella[12] .extended_lut = "off";
defparam \add_sub_cella[12] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[12] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[13] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[12]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[13]~sumout ),
	.cout(\add_sub_cella[13]~COUT ),
	.shareout());
defparam \add_sub_cella[13] .extended_lut = "off";
defparam \add_sub_cella[13] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[13] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[14] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[13]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[14]~sumout ),
	.cout(\add_sub_cella[14]~COUT ),
	.shareout());
defparam \add_sub_cella[14] .extended_lut = "off";
defparam \add_sub_cella[14] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[14] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[15] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[14]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[15]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[15] .extended_lut = "off";
defparam \add_sub_cella[15] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[15] .shared_arith = "off";

endmodule

module nco_test_cordic_zxor_1p_lpm_6 (
	corz_14,
	corz_13,
	corz_12,
	corz_11,
	corz_10,
	corz_9,
	corz_8,
	corz_7,
	corz_6,
	corz_5,
	corz_4,
	corz_3,
	corz_2,
	corz_1,
	corz_0,
	sin_o_0,
	dffe16,
	corx_10,
	dffe15,
	dffe14,
	dffe13,
	dffe12,
	dffe11,
	dffe10,
	dffe9,
	dffe8,
	dffe7,
	dffe6,
	dffe5,
	dffe4,
	dffe3,
	dffe2,
	dffe1,
	dffe161,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	corz_14;
input 	corz_13;
input 	corz_12;
input 	corz_11;
input 	corz_10;
input 	corz_9;
input 	corz_8;
input 	corz_7;
input 	corz_6;
input 	corz_5;
input 	corz_4;
input 	corz_3;
input 	corz_2;
input 	corz_1;
input 	corz_0;
input 	sin_o_0;
output 	dffe16;
input 	corx_10;
output 	dffe15;
output 	dffe14;
output 	dffe13;
output 	dffe12;
output 	dffe11;
output 	dffe10;
output 	dffe9;
output 	dffe8;
output 	dffe7;
output 	dffe6;
output 	dffe5;
output 	dffe4;
output 	dffe3;
output 	dffe2;
output 	dffe1;
output 	dffe161;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[14]~q ;
wire \a[13]~q ;
wire \a[12]~q ;
wire \a[11]~q ;
wire \a[10]~q ;
wire \a[9]~q ;
wire \a[8]~q ;
wire \a[7]~q ;
wire \a[6]~q ;
wire \a[5]~q ;
wire \a[4]~q ;
wire \a[3]~q ;
wire \a[2]~q ;
wire \a[1]~q ;
wire \a[0]~q ;


nco_test_lpm_add_sub_46 u0(
	.a_14(\a[14]~q ),
	.a_13(\a[13]~q ),
	.a_12(\a[12]~q ),
	.a_11(\a[11]~q ),
	.a_10(\a[10]~q ),
	.a_9(\a[9]~q ),
	.a_8(\a[8]~q ),
	.a_7(\a[7]~q ),
	.a_6(\a[6]~q ),
	.a_5(\a[5]~q ),
	.a_4(\a[4]~q ),
	.a_3(\a[3]~q ),
	.a_2(\a[2]~q ),
	.a_1(\a[1]~q ),
	.a_0(\a[0]~q ),
	.dffe16(dffe16),
	.corx_10(corx_10),
	.dffe15(dffe15),
	.dffe14(dffe14),
	.dffe13(dffe13),
	.dffe12(dffe12),
	.dffe11(dffe11),
	.dffe10(dffe10),
	.dffe9(dffe9),
	.dffe8(dffe8),
	.dffe7(dffe7),
	.dffe6(dffe6),
	.dffe5(dffe5),
	.dffe4(dffe4),
	.dffe3(dffe3),
	.dffe2(dffe2),
	.dffe1(dffe1),
	.dffe161(dffe161),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[14] (
	.clk(clk),
	.d(corz_14),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

dffeas \a[13] (
	.clk(clk),
	.d(corz_13),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

dffeas \a[12] (
	.clk(clk),
	.d(corz_12),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

dffeas \a[11] (
	.clk(clk),
	.d(corz_11),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

dffeas \a[10] (
	.clk(clk),
	.d(corz_10),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

dffeas \a[9] (
	.clk(clk),
	.d(corz_9),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

dffeas \a[8] (
	.clk(clk),
	.d(corz_8),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

dffeas \a[7] (
	.clk(clk),
	.d(corz_7),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

dffeas \a[6] (
	.clk(clk),
	.d(corz_6),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

dffeas \a[5] (
	.clk(clk),
	.d(corz_5),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \a[4] (
	.clk(clk),
	.d(corz_4),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \a[3] (
	.clk(clk),
	.d(corz_3),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \a[2] (
	.clk(clk),
	.d(corz_2),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \a[1] (
	.clk(clk),
	.d(corz_1),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \a[0] (
	.clk(clk),
	.d(corz_0),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

endmodule

module nco_test_cordic_zxor_1p_lpm_7 (
	sin_o_0,
	dffe16,
	dffe15,
	dffe14,
	dffe161,
	dffe13,
	dffe12,
	dffe151,
	dffe11,
	dffe141,
	dffe10,
	dffe131,
	dffe9,
	dffe121,
	dffe8,
	dffe111,
	dffe7,
	dffe101,
	dffe6,
	dffe91,
	dffe5,
	dffe81,
	dffe4,
	dffe71,
	dffe3,
	dffe61,
	dffe2,
	dffe51,
	dffe1,
	dffe41,
	dffe31,
	dffe21,
	dffe17,
	dffe162,
	dffe163,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	sin_o_0;
output 	dffe16;
output 	dffe15;
output 	dffe14;
input 	dffe161;
output 	dffe13;
output 	dffe12;
input 	dffe151;
output 	dffe11;
input 	dffe141;
output 	dffe10;
input 	dffe131;
output 	dffe9;
input 	dffe121;
output 	dffe8;
input 	dffe111;
output 	dffe7;
input 	dffe101;
output 	dffe6;
input 	dffe91;
output 	dffe5;
input 	dffe81;
output 	dffe4;
input 	dffe71;
output 	dffe3;
input 	dffe61;
output 	dffe2;
input 	dffe51;
output 	dffe1;
input 	dffe41;
input 	dffe31;
input 	dffe21;
input 	dffe17;
input 	dffe162;
output 	dffe163;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[15]~q ;
wire \xordvalue[0]~q ;
wire \Add0~1_sumout ;
wire \a[14]~q ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \a[13]~q ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \a[12]~q ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \a[11]~q ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \a[10]~q ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \a[9]~q ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \a[8]~q ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \a[7]~q ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \a[6]~q ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \a[5]~q ;
wire \xordvalue[3]~q ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \a[4]~q ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \a[3]~q ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~51 ;
wire \a[2]~q ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~55 ;
wire \a[1]~q ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~59 ;
wire \a[0]~q ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~63 ;


nco_test_lpm_add_sub_42 u0(
	.a_15(\a[15]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_14(\a[14]~q ),
	.a_13(\a[13]~q ),
	.a_12(\a[12]~q ),
	.a_11(\a[11]~q ),
	.a_10(\a[10]~q ),
	.a_9(\a[9]~q ),
	.a_8(\a[8]~q ),
	.a_7(\a[7]~q ),
	.a_6(\a[6]~q ),
	.a_5(\a[5]~q ),
	.xordvalue_3(\xordvalue[3]~q ),
	.a_4(\a[4]~q ),
	.a_3(\a[3]~q ),
	.a_2(\a[2]~q ),
	.a_1(\a[1]~q ),
	.a_0(\a[0]~q ),
	.dffe16(dffe16),
	.dffe15(dffe15),
	.dffe14(dffe14),
	.dffe13(dffe13),
	.dffe12(dffe12),
	.dffe11(dffe11),
	.dffe10(dffe10),
	.dffe9(dffe9),
	.dffe8(dffe8),
	.dffe7(dffe7),
	.dffe6(dffe6),
	.dffe5(dffe5),
	.dffe4(dffe4),
	.dffe3(dffe3),
	.dffe2(dffe2),
	.dffe1(dffe1),
	.dffe161(dffe163),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(dffe161),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "on";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~5 .shared_arith = "on";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~9 .shared_arith = "on";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~13 .shared_arith = "on";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~17 .shared_arith = "on";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "on";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~25 .shared_arith = "on";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~29 .shared_arith = "on";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~33 .shared_arith = "on";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~37 .shared_arith = "on";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

dffeas \xordvalue[3] (
	.clk(clk),
	.d(dffe162),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[3]~q ),
	.prn(vcc));
defparam \xordvalue[3] .is_wysiwyg = "true";
defparam \xordvalue[3] .power_up = "low";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(\Add0~47 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~41 .shared_arith = "on";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(\Add0~51 ),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout(\Add0~47 ));
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~45 .shared_arith = "on";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(\Add0~55 ),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout(\Add0~51 ));
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~49 .shared_arith = "on";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(\Add0~59 ),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout(\Add0~55 ));
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~53 .shared_arith = "on";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(\Add0~63 ),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout(\Add0~59 ));
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~57 .shared_arith = "on";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!dffe17),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout(\Add0~63 ));
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add0~61 .shared_arith = "on";

endmodule

module nco_test_lpm_add_sub_42 (
	a_15,
	xordvalue_0,
	a_14,
	a_13,
	a_12,
	a_11,
	a_10,
	a_9,
	a_8,
	a_7,
	a_6,
	a_5,
	xordvalue_3,
	a_4,
	a_3,
	a_2,
	a_1,
	a_0,
	dffe16,
	dffe15,
	dffe14,
	dffe13,
	dffe12,
	dffe11,
	dffe10,
	dffe9,
	dffe8,
	dffe7,
	dffe6,
	dffe5,
	dffe4,
	dffe3,
	dffe2,
	dffe1,
	dffe161,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_15;
input 	xordvalue_0;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_10;
input 	a_9;
input 	a_8;
input 	a_7;
input 	a_6;
input 	a_5;
input 	xordvalue_3;
input 	a_4;
input 	a_3;
input 	a_2;
input 	a_1;
input 	a_0;
output 	dffe16;
output 	dffe15;
output 	dffe14;
output 	dffe13;
output 	dffe12;
output 	dffe11;
output 	dffe10;
output 	dffe9;
output 	dffe8;
output 	dffe7;
output 	dffe6;
output 	dffe5;
output 	dffe4;
output 	dffe3;
output 	dffe2;
output 	dffe1;
output 	dffe161;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_add_sub_hdg_6 auto_generated(
	.a_15(a_15),
	.xordvalue_0(xordvalue_0),
	.a_14(a_14),
	.a_13(a_13),
	.a_12(a_12),
	.a_11(a_11),
	.a_10(a_10),
	.a_9(a_9),
	.a_8(a_8),
	.a_7(a_7),
	.a_6(a_6),
	.a_5(a_5),
	.xordvalue_3(xordvalue_3),
	.a_4(a_4),
	.a_3(a_3),
	.a_2(a_2),
	.a_1(a_1),
	.a_0(a_0),
	.dffe161(dffe16),
	.dffe151(dffe15),
	.dffe141(dffe14),
	.dffe131(dffe13),
	.dffe121(dffe12),
	.dffe111(dffe11),
	.dffe101(dffe10),
	.dffe91(dffe9),
	.dffe81(dffe8),
	.dffe71(dffe7),
	.dffe61(dffe6),
	.dffe51(dffe5),
	.dffe41(dffe4),
	.dffe31(dffe3),
	.dffe21(dffe2),
	.dffe17(dffe1),
	.dffe162(dffe161),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module nco_test_add_sub_hdg_6 (
	a_15,
	xordvalue_0,
	a_14,
	a_13,
	a_12,
	a_11,
	a_10,
	a_9,
	a_8,
	a_7,
	a_6,
	a_5,
	xordvalue_3,
	a_4,
	a_3,
	a_2,
	a_1,
	a_0,
	dffe161,
	dffe151,
	dffe141,
	dffe131,
	dffe121,
	dffe111,
	dffe101,
	dffe91,
	dffe81,
	dffe71,
	dffe61,
	dffe51,
	dffe41,
	dffe31,
	dffe21,
	dffe17,
	dffe162,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_15;
input 	xordvalue_0;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_10;
input 	a_9;
input 	a_8;
input 	a_7;
input 	a_6;
input 	a_5;
input 	xordvalue_3;
input 	a_4;
input 	a_3;
input 	a_2;
input 	a_1;
input 	a_0;
output 	dffe161;
output 	dffe151;
output 	dffe141;
output 	dffe131;
output 	dffe121;
output 	dffe111;
output 	dffe101;
output 	dffe91;
output 	dffe81;
output 	dffe71;
output 	dffe61;
output 	dffe51;
output 	dffe41;
output 	dffe31;
output 	dffe21;
output 	dffe17;
output 	dffe162;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~COUT ;
wire \add_sub_cella[12]~COUT ;
wire \add_sub_cella[13]~COUT ;
wire \add_sub_cella[14]~COUT ;
wire \add_sub_cella[15]~sumout ;
wire \add_sub_cella[14]~sumout ;
wire \add_sub_cella[13]~sumout ;
wire \add_sub_cella[12]~sumout ;
wire \add_sub_cella[11]~sumout ;
wire \add_sub_cella[10]~sumout ;
wire \add_sub_cella[9]~sumout ;
wire \add_sub_cella[8]~sumout ;
wire \add_sub_cella[7]~sumout ;
wire \add_sub_cella[6]~sumout ;
wire \add_sub_cella[5]~sumout ;
wire \add_sub_cella[4]~sumout ;
wire \add_sub_cella[3]~sumout ;
wire \add_sub_cella[2]~sumout ;
wire \add_sub_cella[1]~sumout ;
wire \add_sub_cella[0]~sumout ;


dffeas dffe16(
	.clk(clock),
	.d(\add_sub_cella[15]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe161),
	.prn(vcc));
defparam dffe16.is_wysiwyg = "true";
defparam dffe16.power_up = "low";

dffeas dffe15(
	.clk(clock),
	.d(\add_sub_cella[14]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe151),
	.prn(vcc));
defparam dffe15.is_wysiwyg = "true";
defparam dffe15.power_up = "low";

dffeas dffe14(
	.clk(clock),
	.d(\add_sub_cella[13]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe141),
	.prn(vcc));
defparam dffe14.is_wysiwyg = "true";
defparam dffe14.power_up = "low";

dffeas dffe13(
	.clk(clock),
	.d(\add_sub_cella[12]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe131),
	.prn(vcc));
defparam dffe13.is_wysiwyg = "true";
defparam dffe13.power_up = "low";

dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe17),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

arriav_lcell_comb \dffe16~_wirecell (
	.dataa(!dffe161),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(dffe162),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffe16~_wirecell .extended_lut = "off";
defparam \dffe16~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dffe16~_wirecell .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_3),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_3),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(\add_sub_cella[11]~COUT ),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[12] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[11]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[12]~sumout ),
	.cout(\add_sub_cella[12]~COUT ),
	.shareout());
defparam \add_sub_cella[12] .extended_lut = "off";
defparam \add_sub_cella[12] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[12] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[13] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[12]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[13]~sumout ),
	.cout(\add_sub_cella[13]~COUT ),
	.shareout());
defparam \add_sub_cella[13] .extended_lut = "off";
defparam \add_sub_cella[13] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[13] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[14] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[13]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[14]~sumout ),
	.cout(\add_sub_cella[14]~COUT ),
	.shareout());
defparam \add_sub_cella[14] .extended_lut = "off";
defparam \add_sub_cella[14] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[14] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[15] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[14]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[15]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[15] .extended_lut = "off";
defparam \add_sub_cella[15] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[15] .shared_arith = "off";

endmodule

module nco_test_cordic_zxor_1p_lpm_8 (
	sin_o_0,
	dffe16,
	dffe15,
	dffe14,
	dffe161,
	dffe13,
	dffe12,
	dffe151,
	dffe11,
	dffe141,
	dffe10,
	dffe131,
	dffe9,
	dffe121,
	dffe8,
	dffe111,
	dffe7,
	dffe101,
	dffe6,
	dffe91,
	dffe5,
	dffe81,
	dffe4,
	dffe71,
	dffe3,
	dffe61,
	dffe2,
	dffe51,
	dffe1,
	dffe41,
	dffe31,
	dffe21,
	dffe17,
	dffe162,
	dffe163,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	sin_o_0;
output 	dffe16;
output 	dffe15;
output 	dffe14;
input 	dffe161;
output 	dffe13;
output 	dffe12;
input 	dffe151;
output 	dffe11;
input 	dffe141;
output 	dffe10;
input 	dffe131;
output 	dffe9;
input 	dffe121;
output 	dffe8;
input 	dffe111;
output 	dffe7;
input 	dffe101;
output 	dffe6;
input 	dffe91;
output 	dffe5;
input 	dffe81;
output 	dffe4;
input 	dffe71;
output 	dffe3;
input 	dffe61;
output 	dffe2;
input 	dffe51;
output 	dffe1;
input 	dffe41;
input 	dffe31;
input 	dffe21;
input 	dffe17;
input 	dffe162;
output 	dffe163;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[15]~q ;
wire \xordvalue[0]~q ;
wire \Add0~1_sumout ;
wire \a[14]~q ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \a[13]~q ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \a[12]~q ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \a[11]~q ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \a[10]~q ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \a[9]~q ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \a[8]~q ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \a[7]~q ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \a[6]~q ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \a[5]~q ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \a[4]~q ;
wire \xordvalue[2]~q ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \a[3]~q ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~51 ;
wire \a[2]~q ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~55 ;
wire \a[1]~q ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~59 ;
wire \a[0]~q ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~63 ;


nco_test_lpm_add_sub_43 u0(
	.a_15(\a[15]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_14(\a[14]~q ),
	.a_13(\a[13]~q ),
	.a_12(\a[12]~q ),
	.a_11(\a[11]~q ),
	.a_10(\a[10]~q ),
	.a_9(\a[9]~q ),
	.a_8(\a[8]~q ),
	.a_7(\a[7]~q ),
	.a_6(\a[6]~q ),
	.a_5(\a[5]~q ),
	.a_4(\a[4]~q ),
	.xordvalue_2(\xordvalue[2]~q ),
	.a_3(\a[3]~q ),
	.a_2(\a[2]~q ),
	.a_1(\a[1]~q ),
	.a_0(\a[0]~q ),
	.dffe16(dffe16),
	.dffe15(dffe15),
	.dffe14(dffe14),
	.dffe13(dffe13),
	.dffe12(dffe12),
	.dffe11(dffe11),
	.dffe10(dffe10),
	.dffe9(dffe9),
	.dffe8(dffe8),
	.dffe7(dffe7),
	.dffe6(dffe6),
	.dffe5(dffe5),
	.dffe4(dffe4),
	.dffe3(dffe3),
	.dffe2(dffe2),
	.dffe1(dffe1),
	.dffe161(dffe163),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(dffe161),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "on";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~5 .shared_arith = "on";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~9 .shared_arith = "on";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~13 .shared_arith = "on";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~17 .shared_arith = "on";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "on";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~25 .shared_arith = "on";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~29 .shared_arith = "on";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~33 .shared_arith = "on";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~37 .shared_arith = "on";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(\Add0~47 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~41 .shared_arith = "on";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

dffeas \xordvalue[2] (
	.clk(clk),
	.d(dffe162),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[2]~q ),
	.prn(vcc));
defparam \xordvalue[2] .is_wysiwyg = "true";
defparam \xordvalue[2] .power_up = "low";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(\Add0~51 ),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout(\Add0~47 ));
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~45 .shared_arith = "on";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(\Add0~55 ),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout(\Add0~51 ));
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~49 .shared_arith = "on";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(\Add0~59 ),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout(\Add0~55 ));
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~53 .shared_arith = "on";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(\Add0~63 ),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout(\Add0~59 ));
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~57 .shared_arith = "on";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!dffe17),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout(\Add0~63 ));
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add0~61 .shared_arith = "on";

endmodule

module nco_test_lpm_add_sub_43 (
	a_15,
	xordvalue_0,
	a_14,
	a_13,
	a_12,
	a_11,
	a_10,
	a_9,
	a_8,
	a_7,
	a_6,
	a_5,
	a_4,
	xordvalue_2,
	a_3,
	a_2,
	a_1,
	a_0,
	dffe16,
	dffe15,
	dffe14,
	dffe13,
	dffe12,
	dffe11,
	dffe10,
	dffe9,
	dffe8,
	dffe7,
	dffe6,
	dffe5,
	dffe4,
	dffe3,
	dffe2,
	dffe1,
	dffe161,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_15;
input 	xordvalue_0;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_10;
input 	a_9;
input 	a_8;
input 	a_7;
input 	a_6;
input 	a_5;
input 	a_4;
input 	xordvalue_2;
input 	a_3;
input 	a_2;
input 	a_1;
input 	a_0;
output 	dffe16;
output 	dffe15;
output 	dffe14;
output 	dffe13;
output 	dffe12;
output 	dffe11;
output 	dffe10;
output 	dffe9;
output 	dffe8;
output 	dffe7;
output 	dffe6;
output 	dffe5;
output 	dffe4;
output 	dffe3;
output 	dffe2;
output 	dffe1;
output 	dffe161;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_add_sub_hdg_7 auto_generated(
	.a_15(a_15),
	.xordvalue_0(xordvalue_0),
	.a_14(a_14),
	.a_13(a_13),
	.a_12(a_12),
	.a_11(a_11),
	.a_10(a_10),
	.a_9(a_9),
	.a_8(a_8),
	.a_7(a_7),
	.a_6(a_6),
	.a_5(a_5),
	.a_4(a_4),
	.xordvalue_2(xordvalue_2),
	.a_3(a_3),
	.a_2(a_2),
	.a_1(a_1),
	.a_0(a_0),
	.dffe161(dffe16),
	.dffe151(dffe15),
	.dffe141(dffe14),
	.dffe131(dffe13),
	.dffe121(dffe12),
	.dffe111(dffe11),
	.dffe101(dffe10),
	.dffe91(dffe9),
	.dffe81(dffe8),
	.dffe71(dffe7),
	.dffe61(dffe6),
	.dffe51(dffe5),
	.dffe41(dffe4),
	.dffe31(dffe3),
	.dffe21(dffe2),
	.dffe17(dffe1),
	.dffe162(dffe161),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module nco_test_add_sub_hdg_7 (
	a_15,
	xordvalue_0,
	a_14,
	a_13,
	a_12,
	a_11,
	a_10,
	a_9,
	a_8,
	a_7,
	a_6,
	a_5,
	a_4,
	xordvalue_2,
	a_3,
	a_2,
	a_1,
	a_0,
	dffe161,
	dffe151,
	dffe141,
	dffe131,
	dffe121,
	dffe111,
	dffe101,
	dffe91,
	dffe81,
	dffe71,
	dffe61,
	dffe51,
	dffe41,
	dffe31,
	dffe21,
	dffe17,
	dffe162,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_15;
input 	xordvalue_0;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_10;
input 	a_9;
input 	a_8;
input 	a_7;
input 	a_6;
input 	a_5;
input 	a_4;
input 	xordvalue_2;
input 	a_3;
input 	a_2;
input 	a_1;
input 	a_0;
output 	dffe161;
output 	dffe151;
output 	dffe141;
output 	dffe131;
output 	dffe121;
output 	dffe111;
output 	dffe101;
output 	dffe91;
output 	dffe81;
output 	dffe71;
output 	dffe61;
output 	dffe51;
output 	dffe41;
output 	dffe31;
output 	dffe21;
output 	dffe17;
output 	dffe162;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~COUT ;
wire \add_sub_cella[12]~COUT ;
wire \add_sub_cella[13]~COUT ;
wire \add_sub_cella[14]~COUT ;
wire \add_sub_cella[15]~sumout ;
wire \add_sub_cella[14]~sumout ;
wire \add_sub_cella[13]~sumout ;
wire \add_sub_cella[12]~sumout ;
wire \add_sub_cella[11]~sumout ;
wire \add_sub_cella[10]~sumout ;
wire \add_sub_cella[9]~sumout ;
wire \add_sub_cella[8]~sumout ;
wire \add_sub_cella[7]~sumout ;
wire \add_sub_cella[6]~sumout ;
wire \add_sub_cella[5]~sumout ;
wire \add_sub_cella[4]~sumout ;
wire \add_sub_cella[3]~sumout ;
wire \add_sub_cella[2]~sumout ;
wire \add_sub_cella[1]~sumout ;
wire \add_sub_cella[0]~sumout ;


dffeas dffe16(
	.clk(clock),
	.d(\add_sub_cella[15]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe161),
	.prn(vcc));
defparam dffe16.is_wysiwyg = "true";
defparam dffe16.power_up = "low";

dffeas dffe15(
	.clk(clock),
	.d(\add_sub_cella[14]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe151),
	.prn(vcc));
defparam dffe15.is_wysiwyg = "true";
defparam dffe15.power_up = "low";

dffeas dffe14(
	.clk(clock),
	.d(\add_sub_cella[13]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe141),
	.prn(vcc));
defparam dffe14.is_wysiwyg = "true";
defparam dffe14.power_up = "low";

dffeas dffe13(
	.clk(clock),
	.d(\add_sub_cella[12]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe131),
	.prn(vcc));
defparam dffe13.is_wysiwyg = "true";
defparam dffe13.power_up = "low";

dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe17),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

arriav_lcell_comb \dffe16~_wirecell (
	.dataa(!dffe161),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(dffe162),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffe16~_wirecell .extended_lut = "off";
defparam \dffe16~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dffe16~_wirecell .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_2),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_2),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(\add_sub_cella[11]~COUT ),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[12] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[11]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[12]~sumout ),
	.cout(\add_sub_cella[12]~COUT ),
	.shareout());
defparam \add_sub_cella[12] .extended_lut = "off";
defparam \add_sub_cella[12] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[12] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[13] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[12]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[13]~sumout ),
	.cout(\add_sub_cella[13]~COUT ),
	.shareout());
defparam \add_sub_cella[13] .extended_lut = "off";
defparam \add_sub_cella[13] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[13] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[14] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[13]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[14]~sumout ),
	.cout(\add_sub_cella[14]~COUT ),
	.shareout());
defparam \add_sub_cella[14] .extended_lut = "off";
defparam \add_sub_cella[14] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[14] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[15] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[14]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[15]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[15] .extended_lut = "off";
defparam \add_sub_cella[15] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[15] .shared_arith = "off";

endmodule

module nco_test_cordic_zxor_1p_lpm_9 (
	sin_o_0,
	dffe16,
	dffe15,
	dffe14,
	dffe161,
	dffe13,
	dffe12,
	dffe151,
	dffe11,
	dffe141,
	dffe10,
	dffe131,
	dffe9,
	dffe121,
	dffe8,
	dffe111,
	dffe7,
	dffe101,
	dffe6,
	dffe91,
	dffe5,
	dffe81,
	dffe4,
	dffe71,
	dffe3,
	dffe61,
	dffe2,
	dffe51,
	dffe1,
	dffe41,
	dffe31,
	dffe21,
	dffe17,
	dffe162,
	dffe163,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	sin_o_0;
output 	dffe16;
output 	dffe15;
output 	dffe14;
input 	dffe161;
output 	dffe13;
output 	dffe12;
input 	dffe151;
output 	dffe11;
input 	dffe141;
output 	dffe10;
input 	dffe131;
output 	dffe9;
input 	dffe121;
output 	dffe8;
input 	dffe111;
output 	dffe7;
input 	dffe101;
output 	dffe6;
input 	dffe91;
output 	dffe5;
input 	dffe81;
output 	dffe4;
input 	dffe71;
output 	dffe3;
input 	dffe61;
output 	dffe2;
input 	dffe51;
output 	dffe1;
input 	dffe41;
input 	dffe31;
input 	dffe21;
input 	dffe17;
input 	dffe162;
output 	dffe163;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[15]~q ;
wire \xordvalue[0]~q ;
wire \Add0~1_sumout ;
wire \a[14]~q ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \a[13]~q ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \a[12]~q ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \a[11]~q ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \a[10]~q ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \a[9]~q ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \a[8]~q ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \a[7]~q ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \a[6]~q ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \a[5]~q ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \a[4]~q ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \a[3]~q ;
wire \xordvalue[1]~q ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~51 ;
wire \a[2]~q ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~55 ;
wire \a[1]~q ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~59 ;
wire \a[0]~q ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~63 ;


nco_test_lpm_add_sub_44 u0(
	.a_15(\a[15]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_14(\a[14]~q ),
	.a_13(\a[13]~q ),
	.a_12(\a[12]~q ),
	.a_11(\a[11]~q ),
	.a_10(\a[10]~q ),
	.a_9(\a[9]~q ),
	.a_8(\a[8]~q ),
	.a_7(\a[7]~q ),
	.a_6(\a[6]~q ),
	.a_5(\a[5]~q ),
	.a_4(\a[4]~q ),
	.a_3(\a[3]~q ),
	.xordvalue_1(\xordvalue[1]~q ),
	.a_2(\a[2]~q ),
	.a_1(\a[1]~q ),
	.a_0(\a[0]~q ),
	.dffe16(dffe16),
	.dffe15(dffe15),
	.dffe14(dffe14),
	.dffe13(dffe13),
	.dffe12(dffe12),
	.dffe11(dffe11),
	.dffe10(dffe10),
	.dffe9(dffe9),
	.dffe8(dffe8),
	.dffe7(dffe7),
	.dffe6(dffe6),
	.dffe5(dffe5),
	.dffe4(dffe4),
	.dffe3(dffe3),
	.dffe2(dffe2),
	.dffe1(dffe1),
	.dffe161(dffe163),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(dffe161),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "on";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~5 .shared_arith = "on";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~9 .shared_arith = "on";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~13 .shared_arith = "on";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~17 .shared_arith = "on";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "on";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~25 .shared_arith = "on";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~29 .shared_arith = "on";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~33 .shared_arith = "on";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~37 .shared_arith = "on";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(\Add0~47 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~41 .shared_arith = "on";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(\Add0~51 ),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout(\Add0~47 ));
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~45 .shared_arith = "on";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

dffeas \xordvalue[1] (
	.clk(clk),
	.d(dffe162),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[1]~q ),
	.prn(vcc));
defparam \xordvalue[1] .is_wysiwyg = "true";
defparam \xordvalue[1] .power_up = "low";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(\Add0~55 ),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout(\Add0~51 ));
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~49 .shared_arith = "on";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(\Add0~59 ),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout(\Add0~55 ));
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~53 .shared_arith = "on";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(\Add0~63 ),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout(\Add0~59 ));
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~57 .shared_arith = "on";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!dffe17),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout(\Add0~63 ));
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add0~61 .shared_arith = "on";

endmodule

module nco_test_lpm_add_sub_44 (
	a_15,
	xordvalue_0,
	a_14,
	a_13,
	a_12,
	a_11,
	a_10,
	a_9,
	a_8,
	a_7,
	a_6,
	a_5,
	a_4,
	a_3,
	xordvalue_1,
	a_2,
	a_1,
	a_0,
	dffe16,
	dffe15,
	dffe14,
	dffe13,
	dffe12,
	dffe11,
	dffe10,
	dffe9,
	dffe8,
	dffe7,
	dffe6,
	dffe5,
	dffe4,
	dffe3,
	dffe2,
	dffe1,
	dffe161,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_15;
input 	xordvalue_0;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_10;
input 	a_9;
input 	a_8;
input 	a_7;
input 	a_6;
input 	a_5;
input 	a_4;
input 	a_3;
input 	xordvalue_1;
input 	a_2;
input 	a_1;
input 	a_0;
output 	dffe16;
output 	dffe15;
output 	dffe14;
output 	dffe13;
output 	dffe12;
output 	dffe11;
output 	dffe10;
output 	dffe9;
output 	dffe8;
output 	dffe7;
output 	dffe6;
output 	dffe5;
output 	dffe4;
output 	dffe3;
output 	dffe2;
output 	dffe1;
output 	dffe161;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_add_sub_hdg_8 auto_generated(
	.a_15(a_15),
	.xordvalue_0(xordvalue_0),
	.a_14(a_14),
	.a_13(a_13),
	.a_12(a_12),
	.a_11(a_11),
	.a_10(a_10),
	.a_9(a_9),
	.a_8(a_8),
	.a_7(a_7),
	.a_6(a_6),
	.a_5(a_5),
	.a_4(a_4),
	.a_3(a_3),
	.xordvalue_1(xordvalue_1),
	.a_2(a_2),
	.a_1(a_1),
	.a_0(a_0),
	.dffe161(dffe16),
	.dffe151(dffe15),
	.dffe141(dffe14),
	.dffe131(dffe13),
	.dffe121(dffe12),
	.dffe111(dffe11),
	.dffe101(dffe10),
	.dffe91(dffe9),
	.dffe81(dffe8),
	.dffe71(dffe7),
	.dffe61(dffe6),
	.dffe51(dffe5),
	.dffe41(dffe4),
	.dffe31(dffe3),
	.dffe21(dffe2),
	.dffe17(dffe1),
	.dffe162(dffe161),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module nco_test_add_sub_hdg_8 (
	a_15,
	xordvalue_0,
	a_14,
	a_13,
	a_12,
	a_11,
	a_10,
	a_9,
	a_8,
	a_7,
	a_6,
	a_5,
	a_4,
	a_3,
	xordvalue_1,
	a_2,
	a_1,
	a_0,
	dffe161,
	dffe151,
	dffe141,
	dffe131,
	dffe121,
	dffe111,
	dffe101,
	dffe91,
	dffe81,
	dffe71,
	dffe61,
	dffe51,
	dffe41,
	dffe31,
	dffe21,
	dffe17,
	dffe162,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_15;
input 	xordvalue_0;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_10;
input 	a_9;
input 	a_8;
input 	a_7;
input 	a_6;
input 	a_5;
input 	a_4;
input 	a_3;
input 	xordvalue_1;
input 	a_2;
input 	a_1;
input 	a_0;
output 	dffe161;
output 	dffe151;
output 	dffe141;
output 	dffe131;
output 	dffe121;
output 	dffe111;
output 	dffe101;
output 	dffe91;
output 	dffe81;
output 	dffe71;
output 	dffe61;
output 	dffe51;
output 	dffe41;
output 	dffe31;
output 	dffe21;
output 	dffe17;
output 	dffe162;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~COUT ;
wire \add_sub_cella[12]~COUT ;
wire \add_sub_cella[13]~COUT ;
wire \add_sub_cella[14]~COUT ;
wire \add_sub_cella[15]~sumout ;
wire \add_sub_cella[14]~sumout ;
wire \add_sub_cella[13]~sumout ;
wire \add_sub_cella[12]~sumout ;
wire \add_sub_cella[11]~sumout ;
wire \add_sub_cella[10]~sumout ;
wire \add_sub_cella[9]~sumout ;
wire \add_sub_cella[8]~sumout ;
wire \add_sub_cella[7]~sumout ;
wire \add_sub_cella[6]~sumout ;
wire \add_sub_cella[5]~sumout ;
wire \add_sub_cella[4]~sumout ;
wire \add_sub_cella[3]~sumout ;
wire \add_sub_cella[2]~sumout ;
wire \add_sub_cella[1]~sumout ;
wire \add_sub_cella[0]~sumout ;


dffeas dffe16(
	.clk(clock),
	.d(\add_sub_cella[15]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe161),
	.prn(vcc));
defparam dffe16.is_wysiwyg = "true";
defparam dffe16.power_up = "low";

dffeas dffe15(
	.clk(clock),
	.d(\add_sub_cella[14]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe151),
	.prn(vcc));
defparam dffe15.is_wysiwyg = "true";
defparam dffe15.power_up = "low";

dffeas dffe14(
	.clk(clock),
	.d(\add_sub_cella[13]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe141),
	.prn(vcc));
defparam dffe14.is_wysiwyg = "true";
defparam dffe14.power_up = "low";

dffeas dffe13(
	.clk(clock),
	.d(\add_sub_cella[12]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe131),
	.prn(vcc));
defparam dffe13.is_wysiwyg = "true";
defparam dffe13.power_up = "low";

dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe17),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

arriav_lcell_comb \dffe16~_wirecell (
	.dataa(!dffe161),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(dffe162),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffe16~_wirecell .extended_lut = "off";
defparam \dffe16~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dffe16~_wirecell .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_1),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_1),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(\add_sub_cella[11]~COUT ),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[12] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[11]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[12]~sumout ),
	.cout(\add_sub_cella[12]~COUT ),
	.shareout());
defparam \add_sub_cella[12] .extended_lut = "off";
defparam \add_sub_cella[12] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[12] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[13] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[12]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[13]~sumout ),
	.cout(\add_sub_cella[13]~COUT ),
	.shareout());
defparam \add_sub_cella[13] .extended_lut = "off";
defparam \add_sub_cella[13] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[13] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[14] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[13]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[14]~sumout ),
	.cout(\add_sub_cella[14]~COUT ),
	.shareout());
defparam \add_sub_cella[14] .extended_lut = "off";
defparam \add_sub_cella[14] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[14] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[15] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[14]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[15]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[15] .extended_lut = "off";
defparam \add_sub_cella[15] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[15] .shared_arith = "off";

endmodule

module nco_test_cordic_zxor_1p_lpm_10 (
	sin_o_0,
	dffe16,
	dffe15,
	dffe14,
	dffe161,
	dffe13,
	dffe12,
	dffe151,
	dffe11,
	dffe141,
	dffe10,
	dffe131,
	dffe9,
	dffe121,
	dffe8,
	dffe111,
	dffe7,
	dffe101,
	dffe6,
	dffe91,
	dffe5,
	dffe81,
	dffe4,
	dffe71,
	dffe3,
	dffe61,
	dffe2,
	dffe51,
	dffe1,
	dffe41,
	dffe31,
	dffe21,
	dffe17,
	dffe162,
	dffe163,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	sin_o_0;
output 	dffe16;
output 	dffe15;
output 	dffe14;
input 	dffe161;
output 	dffe13;
output 	dffe12;
input 	dffe151;
output 	dffe11;
input 	dffe141;
output 	dffe10;
input 	dffe131;
output 	dffe9;
input 	dffe121;
output 	dffe8;
input 	dffe111;
output 	dffe7;
input 	dffe101;
output 	dffe6;
input 	dffe91;
output 	dffe5;
input 	dffe81;
output 	dffe4;
input 	dffe71;
output 	dffe3;
input 	dffe61;
output 	dffe2;
input 	dffe51;
output 	dffe1;
input 	dffe41;
input 	dffe31;
input 	dffe21;
input 	dffe17;
input 	dffe162;
output 	dffe163;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[15]~q ;
wire \xordvalue[10]~q ;
wire \Add0~1_sumout ;
wire \a[14]~q ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \a[13]~q ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \a[12]~q ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \a[11]~q ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \a[10]~q ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \a[9]~q ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \a[8]~q ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \a[7]~q ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \a[6]~q ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \a[5]~q ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \a[4]~q ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \a[3]~q ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~51 ;
wire \a[2]~q ;
wire \xordvalue[0]~q ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~55 ;
wire \a[1]~q ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~59 ;
wire \a[0]~q ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~63 ;


nco_test_lpm_add_sub_45 u0(
	.a_15(\a[15]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.a_14(\a[14]~q ),
	.a_13(\a[13]~q ),
	.a_12(\a[12]~q ),
	.a_11(\a[11]~q ),
	.a_10(\a[10]~q ),
	.a_9(\a[9]~q ),
	.a_8(\a[8]~q ),
	.a_7(\a[7]~q ),
	.a_6(\a[6]~q ),
	.a_5(\a[5]~q ),
	.a_4(\a[4]~q ),
	.a_3(\a[3]~q ),
	.a_2(\a[2]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_1(\a[1]~q ),
	.a_0(\a[0]~q ),
	.dffe16(dffe16),
	.dffe15(dffe15),
	.dffe14(dffe14),
	.dffe13(dffe13),
	.dffe12(dffe12),
	.dffe11(dffe11),
	.dffe10(dffe10),
	.dffe9(dffe9),
	.dffe8(dffe8),
	.dffe7(dffe7),
	.dffe6(dffe6),
	.dffe5(dffe5),
	.dffe4(dffe4),
	.dffe3(dffe3),
	.dffe2(dffe2),
	.dffe1(dffe1),
	.dffe161(dffe163),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(dffe161),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "on";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~5 .shared_arith = "on";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~9 .shared_arith = "on";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~13 .shared_arith = "on";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~17 .shared_arith = "on";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "on";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~25 .shared_arith = "on";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~29 .shared_arith = "on";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~33 .shared_arith = "on";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~37 .shared_arith = "on";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(\Add0~47 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~41 .shared_arith = "on";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(\Add0~51 ),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout(\Add0~47 ));
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~45 .shared_arith = "on";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(\Add0~55 ),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout(\Add0~51 ));
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~49 .shared_arith = "on";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(dffe162),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(\Add0~59 ),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout(\Add0~55 ));
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~53 .shared_arith = "on";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(\Add0~63 ),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout(\Add0~59 ));
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~57 .shared_arith = "on";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!dffe17),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout(\Add0~63 ));
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add0~61 .shared_arith = "on";

endmodule

module nco_test_lpm_add_sub_45 (
	a_15,
	xordvalue_10,
	a_14,
	a_13,
	a_12,
	a_11,
	a_10,
	a_9,
	a_8,
	a_7,
	a_6,
	a_5,
	a_4,
	a_3,
	a_2,
	xordvalue_0,
	a_1,
	a_0,
	dffe16,
	dffe15,
	dffe14,
	dffe13,
	dffe12,
	dffe11,
	dffe10,
	dffe9,
	dffe8,
	dffe7,
	dffe6,
	dffe5,
	dffe4,
	dffe3,
	dffe2,
	dffe1,
	dffe161,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_15;
input 	xordvalue_10;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_10;
input 	a_9;
input 	a_8;
input 	a_7;
input 	a_6;
input 	a_5;
input 	a_4;
input 	a_3;
input 	a_2;
input 	xordvalue_0;
input 	a_1;
input 	a_0;
output 	dffe16;
output 	dffe15;
output 	dffe14;
output 	dffe13;
output 	dffe12;
output 	dffe11;
output 	dffe10;
output 	dffe9;
output 	dffe8;
output 	dffe7;
output 	dffe6;
output 	dffe5;
output 	dffe4;
output 	dffe3;
output 	dffe2;
output 	dffe1;
output 	dffe161;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_add_sub_hdg_9 auto_generated(
	.a_15(a_15),
	.xordvalue_10(xordvalue_10),
	.a_14(a_14),
	.a_13(a_13),
	.a_12(a_12),
	.a_11(a_11),
	.a_10(a_10),
	.a_9(a_9),
	.a_8(a_8),
	.a_7(a_7),
	.a_6(a_6),
	.a_5(a_5),
	.a_4(a_4),
	.a_3(a_3),
	.a_2(a_2),
	.xordvalue_0(xordvalue_0),
	.a_1(a_1),
	.a_0(a_0),
	.dffe161(dffe16),
	.dffe151(dffe15),
	.dffe141(dffe14),
	.dffe131(dffe13),
	.dffe121(dffe12),
	.dffe111(dffe11),
	.dffe101(dffe10),
	.dffe91(dffe9),
	.dffe81(dffe8),
	.dffe71(dffe7),
	.dffe61(dffe6),
	.dffe51(dffe5),
	.dffe41(dffe4),
	.dffe31(dffe3),
	.dffe21(dffe2),
	.dffe17(dffe1),
	.dffe162(dffe161),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module nco_test_add_sub_hdg_9 (
	a_15,
	xordvalue_10,
	a_14,
	a_13,
	a_12,
	a_11,
	a_10,
	a_9,
	a_8,
	a_7,
	a_6,
	a_5,
	a_4,
	a_3,
	a_2,
	xordvalue_0,
	a_1,
	a_0,
	dffe161,
	dffe151,
	dffe141,
	dffe131,
	dffe121,
	dffe111,
	dffe101,
	dffe91,
	dffe81,
	dffe71,
	dffe61,
	dffe51,
	dffe41,
	dffe31,
	dffe21,
	dffe17,
	dffe162,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_15;
input 	xordvalue_10;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_10;
input 	a_9;
input 	a_8;
input 	a_7;
input 	a_6;
input 	a_5;
input 	a_4;
input 	a_3;
input 	a_2;
input 	xordvalue_0;
input 	a_1;
input 	a_0;
output 	dffe161;
output 	dffe151;
output 	dffe141;
output 	dffe131;
output 	dffe121;
output 	dffe111;
output 	dffe101;
output 	dffe91;
output 	dffe81;
output 	dffe71;
output 	dffe61;
output 	dffe51;
output 	dffe41;
output 	dffe31;
output 	dffe21;
output 	dffe17;
output 	dffe162;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~COUT ;
wire \add_sub_cella[12]~COUT ;
wire \add_sub_cella[13]~COUT ;
wire \add_sub_cella[14]~COUT ;
wire \add_sub_cella[15]~sumout ;
wire \add_sub_cella[14]~sumout ;
wire \add_sub_cella[13]~sumout ;
wire \add_sub_cella[12]~sumout ;
wire \add_sub_cella[11]~sumout ;
wire \add_sub_cella[10]~sumout ;
wire \add_sub_cella[9]~sumout ;
wire \add_sub_cella[8]~sumout ;
wire \add_sub_cella[7]~sumout ;
wire \add_sub_cella[6]~sumout ;
wire \add_sub_cella[5]~sumout ;
wire \add_sub_cella[4]~sumout ;
wire \add_sub_cella[3]~sumout ;
wire \add_sub_cella[2]~sumout ;
wire \add_sub_cella[1]~sumout ;
wire \add_sub_cella[0]~sumout ;


dffeas dffe16(
	.clk(clock),
	.d(\add_sub_cella[15]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe161),
	.prn(vcc));
defparam dffe16.is_wysiwyg = "true";
defparam dffe16.power_up = "low";

dffeas dffe15(
	.clk(clock),
	.d(\add_sub_cella[14]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe151),
	.prn(vcc));
defparam dffe15.is_wysiwyg = "true";
defparam dffe15.power_up = "low";

dffeas dffe14(
	.clk(clock),
	.d(\add_sub_cella[13]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe141),
	.prn(vcc));
defparam dffe14.is_wysiwyg = "true";
defparam dffe14.power_up = "low";

dffeas dffe13(
	.clk(clock),
	.d(\add_sub_cella[12]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe131),
	.prn(vcc));
defparam dffe13.is_wysiwyg = "true";
defparam dffe13.power_up = "low";

dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe17),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

arriav_lcell_comb \dffe16~_wirecell (
	.dataa(!dffe161),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(dffe162),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffe16~_wirecell .extended_lut = "off";
defparam \dffe16~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dffe16~_wirecell .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(\add_sub_cella[11]~COUT ),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[12] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[11]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[12]~sumout ),
	.cout(\add_sub_cella[12]~COUT ),
	.shareout());
defparam \add_sub_cella[12] .extended_lut = "off";
defparam \add_sub_cella[12] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[12] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[13] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[12]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[13]~sumout ),
	.cout(\add_sub_cella[13]~COUT ),
	.shareout());
defparam \add_sub_cella[13] .extended_lut = "off";
defparam \add_sub_cella[13] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[13] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[14] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[13]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[14]~sumout ),
	.cout(\add_sub_cella[14]~COUT ),
	.shareout());
defparam \add_sub_cella[14] .extended_lut = "off";
defparam \add_sub_cella[14] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[14] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[15] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[14]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[15]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[15] .extended_lut = "off";
defparam \add_sub_cella[15] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[15] .shared_arith = "off";

endmodule

module nco_test_lpm_add_sub_46 (
	a_14,
	a_13,
	a_12,
	a_11,
	a_10,
	a_9,
	a_8,
	a_7,
	a_6,
	a_5,
	a_4,
	a_3,
	a_2,
	a_1,
	a_0,
	dffe16,
	corx_10,
	dffe15,
	dffe14,
	dffe13,
	dffe12,
	dffe11,
	dffe10,
	dffe9,
	dffe8,
	dffe7,
	dffe6,
	dffe5,
	dffe4,
	dffe3,
	dffe2,
	dffe1,
	dffe161,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_10;
input 	a_9;
input 	a_8;
input 	a_7;
input 	a_6;
input 	a_5;
input 	a_4;
input 	a_3;
input 	a_2;
input 	a_1;
input 	a_0;
output 	dffe16;
input 	corx_10;
output 	dffe15;
output 	dffe14;
output 	dffe13;
output 	dffe12;
output 	dffe11;
output 	dffe10;
output 	dffe9;
output 	dffe8;
output 	dffe7;
output 	dffe6;
output 	dffe5;
output 	dffe4;
output 	dffe3;
output 	dffe2;
output 	dffe1;
output 	dffe161;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_add_sub_hdg_10 auto_generated(
	.a_14(a_14),
	.a_13(a_13),
	.a_12(a_12),
	.a_11(a_11),
	.a_10(a_10),
	.a_9(a_9),
	.a_8(a_8),
	.a_7(a_7),
	.a_6(a_6),
	.a_5(a_5),
	.a_4(a_4),
	.a_3(a_3),
	.a_2(a_2),
	.a_1(a_1),
	.a_0(a_0),
	.dffe161(dffe16),
	.corx_10(corx_10),
	.dffe151(dffe15),
	.dffe141(dffe14),
	.dffe131(dffe13),
	.dffe121(dffe12),
	.dffe111(dffe11),
	.dffe101(dffe10),
	.dffe91(dffe9),
	.dffe81(dffe8),
	.dffe71(dffe7),
	.dffe61(dffe6),
	.dffe51(dffe5),
	.dffe41(dffe4),
	.dffe31(dffe3),
	.dffe21(dffe2),
	.dffe17(dffe1),
	.dffe162(dffe161),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module nco_test_add_sub_hdg_10 (
	a_14,
	a_13,
	a_12,
	a_11,
	a_10,
	a_9,
	a_8,
	a_7,
	a_6,
	a_5,
	a_4,
	a_3,
	a_2,
	a_1,
	a_0,
	dffe161,
	corx_10,
	dffe151,
	dffe141,
	dffe131,
	dffe121,
	dffe111,
	dffe101,
	dffe91,
	dffe81,
	dffe71,
	dffe61,
	dffe51,
	dffe41,
	dffe31,
	dffe21,
	dffe17,
	dffe162,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_10;
input 	a_9;
input 	a_8;
input 	a_7;
input 	a_6;
input 	a_5;
input 	a_4;
input 	a_3;
input 	a_2;
input 	a_1;
input 	a_0;
output 	dffe161;
input 	corx_10;
output 	dffe151;
output 	dffe141;
output 	dffe131;
output 	dffe121;
output 	dffe111;
output 	dffe101;
output 	dffe91;
output 	dffe81;
output 	dffe71;
output 	dffe61;
output 	dffe51;
output 	dffe41;
output 	dffe31;
output 	dffe21;
output 	dffe17;
output 	dffe162;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~COUT ;
wire \add_sub_cella[12]~COUT ;
wire \add_sub_cella[13]~COUT ;
wire \add_sub_cella[14]~COUT ;
wire \add_sub_cella[15]~sumout ;
wire \add_sub_cella[14]~sumout ;
wire \add_sub_cella[13]~sumout ;
wire \add_sub_cella[12]~sumout ;
wire \add_sub_cella[11]~sumout ;
wire \add_sub_cella[10]~sumout ;
wire \add_sub_cella[9]~sumout ;
wire \add_sub_cella[8]~sumout ;
wire \add_sub_cella[7]~sumout ;
wire \add_sub_cella[6]~sumout ;
wire \add_sub_cella[5]~sumout ;
wire \add_sub_cella[4]~sumout ;
wire \add_sub_cella[3]~sumout ;
wire \add_sub_cella[2]~sumout ;
wire \add_sub_cella[1]~sumout ;
wire \add_sub_cella[0]~sumout ;


dffeas dffe16(
	.clk(clock),
	.d(\add_sub_cella[15]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe161),
	.prn(vcc));
defparam dffe16.is_wysiwyg = "true";
defparam dffe16.power_up = "low";

dffeas dffe15(
	.clk(clock),
	.d(\add_sub_cella[14]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe151),
	.prn(vcc));
defparam dffe15.is_wysiwyg = "true";
defparam dffe15.power_up = "low";

dffeas dffe14(
	.clk(clock),
	.d(\add_sub_cella[13]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe141),
	.prn(vcc));
defparam dffe14.is_wysiwyg = "true";
defparam dffe14.power_up = "low";

dffeas dffe13(
	.clk(clock),
	.d(\add_sub_cella[12]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe131),
	.prn(vcc));
defparam dffe13.is_wysiwyg = "true";
defparam dffe13.power_up = "low";

dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe17),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

arriav_lcell_comb \dffe16~_wirecell (
	.dataa(!dffe161),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(dffe162),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffe16~_wirecell .extended_lut = "off";
defparam \dffe16~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dffe16~_wirecell .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h00000000000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h00000000000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h00000000000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h00000000000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h00000000000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h00000000000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h00000000000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h00000000000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h00000000000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h00000000000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h00000000000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(\add_sub_cella[11]~COUT ),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h00000000000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[12] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\add_sub_cella[11]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[12]~sumout ),
	.cout(\add_sub_cella[12]~COUT ),
	.shareout());
defparam \add_sub_cella[12] .extended_lut = "off";
defparam \add_sub_cella[12] .lut_mask = 64'h00000000000000FF;
defparam \add_sub_cella[12] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[13] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\add_sub_cella[12]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[13]~sumout ),
	.cout(\add_sub_cella[13]~COUT ),
	.shareout());
defparam \add_sub_cella[13] .extended_lut = "off";
defparam \add_sub_cella[13] .lut_mask = 64'h00000000000000FF;
defparam \add_sub_cella[13] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[14] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!corx_10),
	.datag(gnd),
	.cin(\add_sub_cella[13]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[14]~sumout ),
	.cout(\add_sub_cella[14]~COUT ),
	.shareout());
defparam \add_sub_cella[14] .extended_lut = "off";
defparam \add_sub_cella[14] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[14] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[15] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\add_sub_cella[14]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[15]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[15] .extended_lut = "off";
defparam \add_sub_cella[15] .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[15] .shared_arith = "off";

endmodule

module nco_test_cordic_zxor_1p_lpm_11 (
	sin_o_0,
	dffe16,
	dffe15,
	dffe14,
	dffe161,
	dffe13,
	dffe12,
	dffe151,
	dffe11,
	dffe141,
	dffe10,
	dffe131,
	dffe9,
	dffe121,
	dffe8,
	dffe111,
	dffe7,
	dffe101,
	dffe6,
	dffe91,
	dffe5,
	dffe81,
	dffe4,
	dffe71,
	dffe3,
	dffe61,
	dffe2,
	dffe51,
	dffe1,
	dffe41,
	dffe31,
	dffe21,
	dffe17,
	dffe162,
	dffe163,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	sin_o_0;
output 	dffe16;
output 	dffe15;
output 	dffe14;
input 	dffe161;
output 	dffe13;
output 	dffe12;
input 	dffe151;
output 	dffe11;
input 	dffe141;
output 	dffe10;
input 	dffe131;
output 	dffe9;
input 	dffe121;
output 	dffe8;
input 	dffe111;
output 	dffe7;
input 	dffe101;
output 	dffe6;
input 	dffe91;
output 	dffe5;
input 	dffe81;
output 	dffe4;
input 	dffe71;
output 	dffe3;
input 	dffe61;
output 	dffe2;
input 	dffe51;
output 	dffe1;
input 	dffe41;
input 	dffe31;
input 	dffe21;
input 	dffe17;
input 	dffe162;
output 	dffe163;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[15]~q ;
wire \xordvalue[0]~q ;
wire \Add0~1_sumout ;
wire \a[14]~q ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \a[13]~q ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \a[12]~q ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \a[11]~q ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \a[10]~q ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \a[9]~q ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \a[8]~q ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \a[7]~q ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \a[6]~q ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \a[5]~q ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \a[4]~q ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \a[3]~q ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~51 ;
wire \a[2]~q ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~55 ;
wire \a[1]~q ;
wire \xordvalue[1]~q ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~59 ;
wire \a[0]~q ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~63 ;


nco_test_lpm_add_sub_47 u0(
	.a_15(\a[15]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_14(\a[14]~q ),
	.a_13(\a[13]~q ),
	.a_12(\a[12]~q ),
	.a_11(\a[11]~q ),
	.a_10(\a[10]~q ),
	.a_9(\a[9]~q ),
	.a_8(\a[8]~q ),
	.a_7(\a[7]~q ),
	.a_6(\a[6]~q ),
	.a_5(\a[5]~q ),
	.a_4(\a[4]~q ),
	.a_3(\a[3]~q ),
	.a_2(\a[2]~q ),
	.a_1(\a[1]~q ),
	.xordvalue_1(\xordvalue[1]~q ),
	.a_0(\a[0]~q ),
	.dffe16(dffe16),
	.dffe15(dffe15),
	.dffe14(dffe14),
	.dffe13(dffe13),
	.dffe12(dffe12),
	.dffe11(dffe11),
	.dffe10(dffe10),
	.dffe9(dffe9),
	.dffe8(dffe8),
	.dffe7(dffe7),
	.dffe6(dffe6),
	.dffe5(dffe5),
	.dffe4(dffe4),
	.dffe3(dffe3),
	.dffe2(dffe2),
	.dffe1(dffe1),
	.dffe161(dffe163),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(dffe161),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "on";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~5 .shared_arith = "on";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~9 .shared_arith = "on";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~13 .shared_arith = "on";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~17 .shared_arith = "on";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "on";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~25 .shared_arith = "on";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~29 .shared_arith = "on";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~33 .shared_arith = "on";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~37 .shared_arith = "on";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(\Add0~47 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~41 .shared_arith = "on";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(\Add0~51 ),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout(\Add0~47 ));
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~45 .shared_arith = "on";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(\Add0~55 ),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout(\Add0~51 ));
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~49 .shared_arith = "on";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(\Add0~59 ),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout(\Add0~55 ));
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~53 .shared_arith = "on";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

dffeas \xordvalue[1] (
	.clk(clk),
	.d(dffe162),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[1]~q ),
	.prn(vcc));
defparam \xordvalue[1] .is_wysiwyg = "true";
defparam \xordvalue[1] .power_up = "low";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(\Add0~63 ),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout(\Add0~59 ));
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~57 .shared_arith = "on";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!dffe17),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout(\Add0~63 ));
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add0~61 .shared_arith = "on";

endmodule

module nco_test_lpm_add_sub_47 (
	a_15,
	xordvalue_0,
	a_14,
	a_13,
	a_12,
	a_11,
	a_10,
	a_9,
	a_8,
	a_7,
	a_6,
	a_5,
	a_4,
	a_3,
	a_2,
	a_1,
	xordvalue_1,
	a_0,
	dffe16,
	dffe15,
	dffe14,
	dffe13,
	dffe12,
	dffe11,
	dffe10,
	dffe9,
	dffe8,
	dffe7,
	dffe6,
	dffe5,
	dffe4,
	dffe3,
	dffe2,
	dffe1,
	dffe161,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_15;
input 	xordvalue_0;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_10;
input 	a_9;
input 	a_8;
input 	a_7;
input 	a_6;
input 	a_5;
input 	a_4;
input 	a_3;
input 	a_2;
input 	a_1;
input 	xordvalue_1;
input 	a_0;
output 	dffe16;
output 	dffe15;
output 	dffe14;
output 	dffe13;
output 	dffe12;
output 	dffe11;
output 	dffe10;
output 	dffe9;
output 	dffe8;
output 	dffe7;
output 	dffe6;
output 	dffe5;
output 	dffe4;
output 	dffe3;
output 	dffe2;
output 	dffe1;
output 	dffe161;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_add_sub_hdg_11 auto_generated(
	.a_15(a_15),
	.xordvalue_0(xordvalue_0),
	.a_14(a_14),
	.a_13(a_13),
	.a_12(a_12),
	.a_11(a_11),
	.a_10(a_10),
	.a_9(a_9),
	.a_8(a_8),
	.a_7(a_7),
	.a_6(a_6),
	.a_5(a_5),
	.a_4(a_4),
	.a_3(a_3),
	.a_2(a_2),
	.a_1(a_1),
	.xordvalue_1(xordvalue_1),
	.a_0(a_0),
	.dffe161(dffe16),
	.dffe151(dffe15),
	.dffe141(dffe14),
	.dffe131(dffe13),
	.dffe121(dffe12),
	.dffe111(dffe11),
	.dffe101(dffe10),
	.dffe91(dffe9),
	.dffe81(dffe8),
	.dffe71(dffe7),
	.dffe61(dffe6),
	.dffe51(dffe5),
	.dffe41(dffe4),
	.dffe31(dffe3),
	.dffe21(dffe2),
	.dffe17(dffe1),
	.dffe162(dffe161),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module nco_test_add_sub_hdg_11 (
	a_15,
	xordvalue_0,
	a_14,
	a_13,
	a_12,
	a_11,
	a_10,
	a_9,
	a_8,
	a_7,
	a_6,
	a_5,
	a_4,
	a_3,
	a_2,
	a_1,
	xordvalue_1,
	a_0,
	dffe161,
	dffe151,
	dffe141,
	dffe131,
	dffe121,
	dffe111,
	dffe101,
	dffe91,
	dffe81,
	dffe71,
	dffe61,
	dffe51,
	dffe41,
	dffe31,
	dffe21,
	dffe17,
	dffe162,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_15;
input 	xordvalue_0;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_10;
input 	a_9;
input 	a_8;
input 	a_7;
input 	a_6;
input 	a_5;
input 	a_4;
input 	a_3;
input 	a_2;
input 	a_1;
input 	xordvalue_1;
input 	a_0;
output 	dffe161;
output 	dffe151;
output 	dffe141;
output 	dffe131;
output 	dffe121;
output 	dffe111;
output 	dffe101;
output 	dffe91;
output 	dffe81;
output 	dffe71;
output 	dffe61;
output 	dffe51;
output 	dffe41;
output 	dffe31;
output 	dffe21;
output 	dffe17;
output 	dffe162;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~COUT ;
wire \add_sub_cella[12]~COUT ;
wire \add_sub_cella[13]~COUT ;
wire \add_sub_cella[14]~COUT ;
wire \add_sub_cella[15]~sumout ;
wire \add_sub_cella[14]~sumout ;
wire \add_sub_cella[13]~sumout ;
wire \add_sub_cella[12]~sumout ;
wire \add_sub_cella[11]~sumout ;
wire \add_sub_cella[10]~sumout ;
wire \add_sub_cella[9]~sumout ;
wire \add_sub_cella[8]~sumout ;
wire \add_sub_cella[7]~sumout ;
wire \add_sub_cella[6]~sumout ;
wire \add_sub_cella[5]~sumout ;
wire \add_sub_cella[4]~sumout ;
wire \add_sub_cella[3]~sumout ;
wire \add_sub_cella[2]~sumout ;
wire \add_sub_cella[1]~sumout ;
wire \add_sub_cella[0]~sumout ;


dffeas dffe16(
	.clk(clock),
	.d(\add_sub_cella[15]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe161),
	.prn(vcc));
defparam dffe16.is_wysiwyg = "true";
defparam dffe16.power_up = "low";

dffeas dffe15(
	.clk(clock),
	.d(\add_sub_cella[14]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe151),
	.prn(vcc));
defparam dffe15.is_wysiwyg = "true";
defparam dffe15.power_up = "low";

dffeas dffe14(
	.clk(clock),
	.d(\add_sub_cella[13]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe141),
	.prn(vcc));
defparam dffe14.is_wysiwyg = "true";
defparam dffe14.power_up = "low";

dffeas dffe13(
	.clk(clock),
	.d(\add_sub_cella[12]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe131),
	.prn(vcc));
defparam dffe13.is_wysiwyg = "true";
defparam dffe13.power_up = "low";

dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe17),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

arriav_lcell_comb \dffe16~_wirecell (
	.dataa(!dffe161),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(dffe162),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffe16~_wirecell .extended_lut = "off";
defparam \dffe16~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dffe16~_wirecell .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_1),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(\add_sub_cella[11]~COUT ),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[12] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[11]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[12]~sumout ),
	.cout(\add_sub_cella[12]~COUT ),
	.shareout());
defparam \add_sub_cella[12] .extended_lut = "off";
defparam \add_sub_cella[12] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[12] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[13] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[12]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[13]~sumout ),
	.cout(\add_sub_cella[13]~COUT ),
	.shareout());
defparam \add_sub_cella[13] .extended_lut = "off";
defparam \add_sub_cella[13] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[13] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[14] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[13]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[14]~sumout ),
	.cout(\add_sub_cella[14]~COUT ),
	.shareout());
defparam \add_sub_cella[14] .extended_lut = "off";
defparam \add_sub_cella[14] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[14] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[15] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[14]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[15]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[15] .extended_lut = "off";
defparam \add_sub_cella[15] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[15] .shared_arith = "off";

endmodule

module nco_test_cordic_zxor_1p_lpm_12 (
	sin_o_0,
	dffe16,
	dffe15,
	dffe14,
	dffe161,
	dffe13,
	dffe12,
	dffe151,
	dffe11,
	dffe141,
	dffe10,
	dffe131,
	dffe9,
	dffe121,
	dffe8,
	dffe111,
	dffe7,
	dffe101,
	dffe6,
	dffe91,
	dffe5,
	dffe81,
	dffe4,
	dffe71,
	dffe3,
	dffe61,
	dffe2,
	dffe51,
	dffe1,
	dffe41,
	dffe31,
	dffe21,
	dffe17,
	dffe162,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	sin_o_0;
output 	dffe16;
output 	dffe15;
output 	dffe14;
input 	dffe161;
output 	dffe13;
output 	dffe12;
input 	dffe151;
output 	dffe11;
input 	dffe141;
output 	dffe10;
input 	dffe131;
output 	dffe9;
input 	dffe121;
output 	dffe8;
input 	dffe111;
output 	dffe7;
input 	dffe101;
output 	dffe6;
input 	dffe91;
output 	dffe5;
input 	dffe81;
output 	dffe4;
input 	dffe71;
output 	dffe3;
input 	dffe61;
output 	dffe2;
input 	dffe51;
output 	dffe1;
input 	dffe41;
input 	dffe31;
input 	dffe21;
input 	dffe17;
input 	dffe162;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[15]~q ;
wire \xordvalue[10]~q ;
wire \Add0~1_sumout ;
wire \a[14]~q ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \a[13]~q ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \a[12]~q ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \a[11]~q ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \a[10]~q ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \a[9]~q ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \a[8]~q ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \a[7]~q ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \a[6]~q ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \a[5]~q ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \a[4]~q ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \a[3]~q ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~51 ;
wire \a[2]~q ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~55 ;
wire \a[1]~q ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~59 ;
wire \a[0]~q ;
wire \xordvalue[0]~q ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~63 ;


nco_test_lpm_add_sub_48 u0(
	.a_15(\a[15]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.a_14(\a[14]~q ),
	.a_13(\a[13]~q ),
	.a_12(\a[12]~q ),
	.a_11(\a[11]~q ),
	.a_10(\a[10]~q ),
	.a_9(\a[9]~q ),
	.a_8(\a[8]~q ),
	.a_7(\a[7]~q ),
	.a_6(\a[6]~q ),
	.a_5(\a[5]~q ),
	.a_4(\a[4]~q ),
	.a_3(\a[3]~q ),
	.a_2(\a[2]~q ),
	.a_1(\a[1]~q ),
	.a_0(\a[0]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.dffe16(dffe16),
	.dffe15(dffe15),
	.dffe14(dffe14),
	.dffe13(dffe13),
	.dffe12(dffe12),
	.dffe11(dffe11),
	.dffe10(dffe10),
	.dffe9(dffe9),
	.dffe8(dffe8),
	.dffe7(dffe7),
	.dffe6(dffe6),
	.dffe5(dffe5),
	.dffe4(dffe4),
	.dffe3(dffe3),
	.dffe2(dffe2),
	.dffe1(dffe1),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(dffe161),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "on";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~5 .shared_arith = "on";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~9 .shared_arith = "on";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~13 .shared_arith = "on";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~17 .shared_arith = "on";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "on";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~25 .shared_arith = "on";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~29 .shared_arith = "on";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~33 .shared_arith = "on";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~37 .shared_arith = "on";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(\Add0~47 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~41 .shared_arith = "on";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(\Add0~51 ),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout(\Add0~47 ));
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~45 .shared_arith = "on";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(\Add0~55 ),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout(\Add0~51 ));
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~49 .shared_arith = "on";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(\Add0~59 ),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout(\Add0~55 ));
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~53 .shared_arith = "on";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(\Add0~63 ),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout(\Add0~59 ));
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~57 .shared_arith = "on";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(dffe162),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!dffe17),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout(\Add0~63 ));
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add0~61 .shared_arith = "on";

endmodule

module nco_test_lpm_add_sub_48 (
	a_15,
	xordvalue_10,
	a_14,
	a_13,
	a_12,
	a_11,
	a_10,
	a_9,
	a_8,
	a_7,
	a_6,
	a_5,
	a_4,
	a_3,
	a_2,
	a_1,
	a_0,
	xordvalue_0,
	dffe16,
	dffe15,
	dffe14,
	dffe13,
	dffe12,
	dffe11,
	dffe10,
	dffe9,
	dffe8,
	dffe7,
	dffe6,
	dffe5,
	dffe4,
	dffe3,
	dffe2,
	dffe1,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_15;
input 	xordvalue_10;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_10;
input 	a_9;
input 	a_8;
input 	a_7;
input 	a_6;
input 	a_5;
input 	a_4;
input 	a_3;
input 	a_2;
input 	a_1;
input 	a_0;
input 	xordvalue_0;
output 	dffe16;
output 	dffe15;
output 	dffe14;
output 	dffe13;
output 	dffe12;
output 	dffe11;
output 	dffe10;
output 	dffe9;
output 	dffe8;
output 	dffe7;
output 	dffe6;
output 	dffe5;
output 	dffe4;
output 	dffe3;
output 	dffe2;
output 	dffe1;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_add_sub_hdg_12 auto_generated(
	.a_15(a_15),
	.xordvalue_10(xordvalue_10),
	.a_14(a_14),
	.a_13(a_13),
	.a_12(a_12),
	.a_11(a_11),
	.a_10(a_10),
	.a_9(a_9),
	.a_8(a_8),
	.a_7(a_7),
	.a_6(a_6),
	.a_5(a_5),
	.a_4(a_4),
	.a_3(a_3),
	.a_2(a_2),
	.a_1(a_1),
	.a_0(a_0),
	.xordvalue_0(xordvalue_0),
	.dffe161(dffe16),
	.dffe151(dffe15),
	.dffe141(dffe14),
	.dffe131(dffe13),
	.dffe121(dffe12),
	.dffe111(dffe11),
	.dffe101(dffe10),
	.dffe91(dffe9),
	.dffe81(dffe8),
	.dffe71(dffe7),
	.dffe61(dffe6),
	.dffe51(dffe5),
	.dffe41(dffe4),
	.dffe31(dffe3),
	.dffe21(dffe2),
	.dffe17(dffe1),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module nco_test_add_sub_hdg_12 (
	a_15,
	xordvalue_10,
	a_14,
	a_13,
	a_12,
	a_11,
	a_10,
	a_9,
	a_8,
	a_7,
	a_6,
	a_5,
	a_4,
	a_3,
	a_2,
	a_1,
	a_0,
	xordvalue_0,
	dffe161,
	dffe151,
	dffe141,
	dffe131,
	dffe121,
	dffe111,
	dffe101,
	dffe91,
	dffe81,
	dffe71,
	dffe61,
	dffe51,
	dffe41,
	dffe31,
	dffe21,
	dffe17,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_15;
input 	xordvalue_10;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_10;
input 	a_9;
input 	a_8;
input 	a_7;
input 	a_6;
input 	a_5;
input 	a_4;
input 	a_3;
input 	a_2;
input 	a_1;
input 	a_0;
input 	xordvalue_0;
output 	dffe161;
output 	dffe151;
output 	dffe141;
output 	dffe131;
output 	dffe121;
output 	dffe111;
output 	dffe101;
output 	dffe91;
output 	dffe81;
output 	dffe71;
output 	dffe61;
output 	dffe51;
output 	dffe41;
output 	dffe31;
output 	dffe21;
output 	dffe17;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~COUT ;
wire \add_sub_cella[12]~COUT ;
wire \add_sub_cella[13]~COUT ;
wire \add_sub_cella[14]~COUT ;
wire \add_sub_cella[15]~sumout ;
wire \add_sub_cella[14]~sumout ;
wire \add_sub_cella[13]~sumout ;
wire \add_sub_cella[12]~sumout ;
wire \add_sub_cella[11]~sumout ;
wire \add_sub_cella[10]~sumout ;
wire \add_sub_cella[9]~sumout ;
wire \add_sub_cella[8]~sumout ;
wire \add_sub_cella[7]~sumout ;
wire \add_sub_cella[6]~sumout ;
wire \add_sub_cella[5]~sumout ;
wire \add_sub_cella[4]~sumout ;
wire \add_sub_cella[3]~sumout ;
wire \add_sub_cella[2]~sumout ;
wire \add_sub_cella[1]~sumout ;
wire \add_sub_cella[0]~sumout ;


dffeas dffe16(
	.clk(clock),
	.d(\add_sub_cella[15]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe161),
	.prn(vcc));
defparam dffe16.is_wysiwyg = "true";
defparam dffe16.power_up = "low";

dffeas dffe15(
	.clk(clock),
	.d(\add_sub_cella[14]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe151),
	.prn(vcc));
defparam dffe15.is_wysiwyg = "true";
defparam dffe15.power_up = "low";

dffeas dffe14(
	.clk(clock),
	.d(\add_sub_cella[13]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe141),
	.prn(vcc));
defparam dffe14.is_wysiwyg = "true";
defparam dffe14.power_up = "low";

dffeas dffe13(
	.clk(clock),
	.d(\add_sub_cella[12]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe131),
	.prn(vcc));
defparam dffe13.is_wysiwyg = "true";
defparam dffe13.power_up = "low";

dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe17),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

arriav_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(\add_sub_cella[11]~COUT ),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[12] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[11]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[12]~sumout ),
	.cout(\add_sub_cella[12]~COUT ),
	.shareout());
defparam \add_sub_cella[12] .extended_lut = "off";
defparam \add_sub_cella[12] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[12] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[13] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[12]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[13]~sumout ),
	.cout(\add_sub_cella[13]~COUT ),
	.shareout());
defparam \add_sub_cella[13] .extended_lut = "off";
defparam \add_sub_cella[13] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[13] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[14] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[13]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[14]~sumout ),
	.cout(\add_sub_cella[14]~COUT ),
	.shareout());
defparam \add_sub_cella[14] .extended_lut = "off";
defparam \add_sub_cella[14] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[14] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[15] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[14]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[15]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[15] .extended_lut = "off";
defparam \add_sub_cella[15] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[15] .shared_arith = "off";

endmodule

module nco_test_cordic_zxor_1p_lpm_13 (
	sin_o_0,
	dffe16,
	dffe15,
	dffe14,
	dffe161,
	dffe13,
	dffe12,
	dffe151,
	dffe11,
	dffe141,
	dffe10,
	dffe131,
	dffe9,
	dffe121,
	dffe8,
	dffe111,
	dffe7,
	dffe101,
	dffe6,
	dffe91,
	dffe5,
	dffe81,
	dffe4,
	dffe71,
	dffe3,
	dffe61,
	dffe2,
	dffe51,
	dffe1,
	dffe41,
	dffe31,
	dffe21,
	dffe17,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	sin_o_0;
output 	dffe16;
output 	dffe15;
output 	dffe14;
input 	dffe161;
output 	dffe13;
output 	dffe12;
input 	dffe151;
output 	dffe11;
input 	dffe141;
output 	dffe10;
input 	dffe131;
output 	dffe9;
input 	dffe121;
output 	dffe8;
input 	dffe111;
output 	dffe7;
input 	dffe101;
output 	dffe6;
input 	dffe91;
output 	dffe5;
input 	dffe81;
output 	dffe4;
input 	dffe71;
output 	dffe3;
input 	dffe61;
output 	dffe2;
input 	dffe51;
output 	dffe1;
input 	dffe41;
input 	dffe31;
input 	dffe21;
input 	dffe17;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[15]~q ;
wire \xordvalue[0]~q ;
wire \Add0~1_sumout ;
wire \a[14]~q ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \a[13]~q ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \a[12]~q ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \a[11]~q ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \a[10]~q ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \a[9]~q ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \a[8]~q ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \a[7]~q ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \a[6]~q ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \a[5]~q ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \a[4]~q ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \a[3]~q ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~51 ;
wire \a[2]~q ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~55 ;
wire \a[1]~q ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~59 ;
wire \a[0]~q ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~63 ;


nco_test_lpm_add_sub_49 u0(
	.a_15(\a[15]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_14(\a[14]~q ),
	.a_13(\a[13]~q ),
	.a_12(\a[12]~q ),
	.a_11(\a[11]~q ),
	.a_10(\a[10]~q ),
	.a_9(\a[9]~q ),
	.a_8(\a[8]~q ),
	.a_7(\a[7]~q ),
	.a_6(\a[6]~q ),
	.a_5(\a[5]~q ),
	.a_4(\a[4]~q ),
	.a_3(\a[3]~q ),
	.a_2(\a[2]~q ),
	.a_1(\a[1]~q ),
	.a_0(\a[0]~q ),
	.dffe16(dffe16),
	.dffe15(dffe15),
	.dffe14(dffe14),
	.dffe13(dffe13),
	.dffe12(dffe12),
	.dffe11(dffe11),
	.dffe10(dffe10),
	.dffe9(dffe9),
	.dffe8(dffe8),
	.dffe7(dffe7),
	.dffe6(dffe6),
	.dffe5(dffe5),
	.dffe4(dffe4),
	.dffe3(dffe3),
	.dffe2(dffe2),
	.dffe1(dffe1),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(dffe161),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "on";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~5 .shared_arith = "on";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~9 .shared_arith = "on";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~13 .shared_arith = "on";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~17 .shared_arith = "on";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "on";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~25 .shared_arith = "on";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~29 .shared_arith = "on";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~33 .shared_arith = "on";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~37 .shared_arith = "on";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(\Add0~47 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~41 .shared_arith = "on";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(\Add0~51 ),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout(\Add0~47 ));
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~45 .shared_arith = "on";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(\Add0~55 ),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout(\Add0~51 ));
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~49 .shared_arith = "on";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(\Add0~59 ),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout(\Add0~55 ));
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~53 .shared_arith = "on";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(\Add0~63 ),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout(\Add0~59 ));
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~57 .shared_arith = "on";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!dffe17),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout(\Add0~63 ));
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add0~61 .shared_arith = "on";

endmodule

module nco_test_lpm_add_sub_49 (
	a_15,
	xordvalue_0,
	a_14,
	a_13,
	a_12,
	a_11,
	a_10,
	a_9,
	a_8,
	a_7,
	a_6,
	a_5,
	a_4,
	a_3,
	a_2,
	a_1,
	a_0,
	dffe16,
	dffe15,
	dffe14,
	dffe13,
	dffe12,
	dffe11,
	dffe10,
	dffe9,
	dffe8,
	dffe7,
	dffe6,
	dffe5,
	dffe4,
	dffe3,
	dffe2,
	dffe1,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_15;
input 	xordvalue_0;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_10;
input 	a_9;
input 	a_8;
input 	a_7;
input 	a_6;
input 	a_5;
input 	a_4;
input 	a_3;
input 	a_2;
input 	a_1;
input 	a_0;
output 	dffe16;
output 	dffe15;
output 	dffe14;
output 	dffe13;
output 	dffe12;
output 	dffe11;
output 	dffe10;
output 	dffe9;
output 	dffe8;
output 	dffe7;
output 	dffe6;
output 	dffe5;
output 	dffe4;
output 	dffe3;
output 	dffe2;
output 	dffe1;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_add_sub_hdg_13 auto_generated(
	.a_15(a_15),
	.xordvalue_0(xordvalue_0),
	.a_14(a_14),
	.a_13(a_13),
	.a_12(a_12),
	.a_11(a_11),
	.a_10(a_10),
	.a_9(a_9),
	.a_8(a_8),
	.a_7(a_7),
	.a_6(a_6),
	.a_5(a_5),
	.a_4(a_4),
	.a_3(a_3),
	.a_2(a_2),
	.a_1(a_1),
	.a_0(a_0),
	.dffe161(dffe16),
	.dffe151(dffe15),
	.dffe141(dffe14),
	.dffe131(dffe13),
	.dffe121(dffe12),
	.dffe111(dffe11),
	.dffe101(dffe10),
	.dffe91(dffe9),
	.dffe81(dffe8),
	.dffe71(dffe7),
	.dffe61(dffe6),
	.dffe51(dffe5),
	.dffe41(dffe4),
	.dffe31(dffe3),
	.dffe21(dffe2),
	.dffe17(dffe1),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module nco_test_add_sub_hdg_13 (
	a_15,
	xordvalue_0,
	a_14,
	a_13,
	a_12,
	a_11,
	a_10,
	a_9,
	a_8,
	a_7,
	a_6,
	a_5,
	a_4,
	a_3,
	a_2,
	a_1,
	a_0,
	dffe161,
	dffe151,
	dffe141,
	dffe131,
	dffe121,
	dffe111,
	dffe101,
	dffe91,
	dffe81,
	dffe71,
	dffe61,
	dffe51,
	dffe41,
	dffe31,
	dffe21,
	dffe17,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_15;
input 	xordvalue_0;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_10;
input 	a_9;
input 	a_8;
input 	a_7;
input 	a_6;
input 	a_5;
input 	a_4;
input 	a_3;
input 	a_2;
input 	a_1;
input 	a_0;
output 	dffe161;
output 	dffe151;
output 	dffe141;
output 	dffe131;
output 	dffe121;
output 	dffe111;
output 	dffe101;
output 	dffe91;
output 	dffe81;
output 	dffe71;
output 	dffe61;
output 	dffe51;
output 	dffe41;
output 	dffe31;
output 	dffe21;
output 	dffe17;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~COUT ;
wire \add_sub_cella[12]~COUT ;
wire \add_sub_cella[13]~COUT ;
wire \add_sub_cella[14]~COUT ;
wire \add_sub_cella[15]~sumout ;
wire \add_sub_cella[14]~sumout ;
wire \add_sub_cella[13]~sumout ;
wire \add_sub_cella[12]~sumout ;
wire \add_sub_cella[11]~sumout ;
wire \add_sub_cella[10]~sumout ;
wire \add_sub_cella[9]~sumout ;
wire \add_sub_cella[8]~sumout ;
wire \add_sub_cella[7]~sumout ;
wire \add_sub_cella[6]~sumout ;
wire \add_sub_cella[5]~sumout ;
wire \add_sub_cella[4]~sumout ;
wire \add_sub_cella[3]~sumout ;
wire \add_sub_cella[2]~sumout ;
wire \add_sub_cella[1]~sumout ;
wire \add_sub_cella[0]~sumout ;


dffeas dffe16(
	.clk(clock),
	.d(\add_sub_cella[15]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe161),
	.prn(vcc));
defparam dffe16.is_wysiwyg = "true";
defparam dffe16.power_up = "low";

dffeas dffe15(
	.clk(clock),
	.d(\add_sub_cella[14]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe151),
	.prn(vcc));
defparam dffe15.is_wysiwyg = "true";
defparam dffe15.power_up = "low";

dffeas dffe14(
	.clk(clock),
	.d(\add_sub_cella[13]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe141),
	.prn(vcc));
defparam dffe14.is_wysiwyg = "true";
defparam dffe14.power_up = "low";

dffeas dffe13(
	.clk(clock),
	.d(\add_sub_cella[12]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe131),
	.prn(vcc));
defparam dffe13.is_wysiwyg = "true";
defparam dffe13.power_up = "low";

dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe17),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

arriav_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(\add_sub_cella[11]~COUT ),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[12] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[11]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[12]~sumout ),
	.cout(\add_sub_cella[12]~COUT ),
	.shareout());
defparam \add_sub_cella[12] .extended_lut = "off";
defparam \add_sub_cella[12] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[12] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[13] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[12]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[13]~sumout ),
	.cout(\add_sub_cella[13]~COUT ),
	.shareout());
defparam \add_sub_cella[13] .extended_lut = "off";
defparam \add_sub_cella[13] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[13] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[14] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[13]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[14]~sumout ),
	.cout(\add_sub_cella[14]~COUT ),
	.shareout());
defparam \add_sub_cella[14] .extended_lut = "off";
defparam \add_sub_cella[14] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[14] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[15] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[14]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[15]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[15] .extended_lut = "off";
defparam \add_sub_cella[15] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[15] .shared_arith = "off";

endmodule

module nco_test_cordic_zxor_1p_lpm_14 (
	sin_o_0,
	dffe16,
	dffe161,
	dffe15,
	dffe14,
	dffe13,
	dffe12,
	dffe11,
	dffe10,
	dffe9,
	dffe8,
	dffe7,
	dffe6,
	dffe5,
	dffe4,
	dffe3,
	dffe2,
	dffe1,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	sin_o_0;
output 	dffe16;
input 	dffe161;
input 	dffe15;
input 	dffe14;
input 	dffe13;
input 	dffe12;
input 	dffe11;
input 	dffe10;
input 	dffe9;
input 	dffe8;
input 	dffe7;
input 	dffe6;
input 	dffe5;
input 	dffe4;
input 	dffe3;
input 	dffe2;
input 	dffe1;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[15]~q ;
wire \xordvalue[0]~q ;
wire \Add0~1_sumout ;
wire \a[14]~q ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \a[13]~q ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \a[12]~q ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \a[11]~q ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \a[10]~q ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \a[9]~q ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \a[8]~q ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \a[7]~q ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \a[6]~q ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \a[5]~q ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \a[4]~q ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \a[3]~q ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~51 ;
wire \a[2]~q ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~55 ;
wire \a[1]~q ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~59 ;
wire \a[0]~q ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~63 ;


nco_test_lpm_add_sub_50 u0(
	.a_15(\a[15]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_14(\a[14]~q ),
	.a_13(\a[13]~q ),
	.a_12(\a[12]~q ),
	.a_11(\a[11]~q ),
	.a_10(\a[10]~q ),
	.a_9(\a[9]~q ),
	.a_8(\a[8]~q ),
	.a_7(\a[7]~q ),
	.a_6(\a[6]~q ),
	.a_5(\a[5]~q ),
	.a_4(\a[4]~q ),
	.a_3(\a[3]~q ),
	.a_2(\a[2]~q ),
	.a_1(\a[1]~q ),
	.a_0(\a[0]~q ),
	.dffe16(dffe16),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(dffe161),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "on";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe15),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~5 .shared_arith = "on";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe14),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~9 .shared_arith = "on";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe13),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~13 .shared_arith = "on";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe12),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~17 .shared_arith = "on";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe11),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "on";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe10),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~25 .shared_arith = "on";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe9),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~29 .shared_arith = "on";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe8),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~33 .shared_arith = "on";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe7),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~37 .shared_arith = "on";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe6),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(\Add0~47 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~41 .shared_arith = "on";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe5),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(\Add0~51 ),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout(\Add0~47 ));
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~45 .shared_arith = "on";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe4),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(\Add0~55 ),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout(\Add0~51 ));
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~49 .shared_arith = "on";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe3),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(\Add0~59 ),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout(\Add0~55 ));
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~53 .shared_arith = "on";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe2),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(\Add0~63 ),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout(\Add0~59 ));
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~57 .shared_arith = "on";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!dffe1),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout(\Add0~63 ));
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add0~61 .shared_arith = "on";

endmodule

module nco_test_lpm_add_sub_50 (
	a_15,
	xordvalue_0,
	a_14,
	a_13,
	a_12,
	a_11,
	a_10,
	a_9,
	a_8,
	a_7,
	a_6,
	a_5,
	a_4,
	a_3,
	a_2,
	a_1,
	a_0,
	dffe16,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_15;
input 	xordvalue_0;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_10;
input 	a_9;
input 	a_8;
input 	a_7;
input 	a_6;
input 	a_5;
input 	a_4;
input 	a_3;
input 	a_2;
input 	a_1;
input 	a_0;
output 	dffe16;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_add_sub_hdg_14 auto_generated(
	.a_15(a_15),
	.xordvalue_0(xordvalue_0),
	.a_14(a_14),
	.a_13(a_13),
	.a_12(a_12),
	.a_11(a_11),
	.a_10(a_10),
	.a_9(a_9),
	.a_8(a_8),
	.a_7(a_7),
	.a_6(a_6),
	.a_5(a_5),
	.a_4(a_4),
	.a_3(a_3),
	.a_2(a_2),
	.a_1(a_1),
	.a_0(a_0),
	.dffe161(dffe16),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module nco_test_add_sub_hdg_14 (
	a_15,
	xordvalue_0,
	a_14,
	a_13,
	a_12,
	a_11,
	a_10,
	a_9,
	a_8,
	a_7,
	a_6,
	a_5,
	a_4,
	a_3,
	a_2,
	a_1,
	a_0,
	dffe161,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_15;
input 	xordvalue_0;
input 	a_14;
input 	a_13;
input 	a_12;
input 	a_11;
input 	a_10;
input 	a_9;
input 	a_8;
input 	a_7;
input 	a_6;
input 	a_5;
input 	a_4;
input 	a_3;
input 	a_2;
input 	a_1;
input 	a_0;
output 	dffe161;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~COUT ;
wire \add_sub_cella[12]~COUT ;
wire \add_sub_cella[13]~COUT ;
wire \add_sub_cella[14]~COUT ;
wire \add_sub_cella[15]~sumout ;


dffeas dffe16(
	.clk(clock),
	.d(\add_sub_cella[15]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe161),
	.prn(vcc));
defparam dffe16.is_wysiwyg = "true";
defparam dffe16.power_up = "low";

arriav_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[11]~COUT ),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[12] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[11]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[12]~COUT ),
	.shareout());
defparam \add_sub_cella[12] .extended_lut = "off";
defparam \add_sub_cella[12] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[12] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[13] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[12]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[13]~COUT ),
	.shareout());
defparam \add_sub_cella[13] .extended_lut = "off";
defparam \add_sub_cella[13] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[13] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[14] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[13]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[14]~COUT ),
	.shareout());
defparam \add_sub_cella[14] .extended_lut = "off";
defparam \add_sub_cella[14] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[14] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[15] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[14]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[15]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[15] .extended_lut = "off";
defparam \add_sub_cella[15] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[15] .shared_arith = "off";

endmodule

module nco_test_cordic_zxor_1p_lpm_15 (
	a_0,
	sin_o_0,
	dffe16,
	dffe15,
	dffe161,
	dffe14,
	dffe13,
	dffe12,
	dffe151,
	dffe11,
	dffe141,
	dffe10,
	dffe131,
	dffe9,
	dffe121,
	dffe8,
	dffe111,
	dffe7,
	dffe101,
	dffe6,
	dffe91,
	dffe5,
	dffe81,
	dffe4,
	dffe71,
	dffe3,
	dffe61,
	dffe2,
	dffe51,
	dffe1,
	dffe41,
	dffe31,
	dffe21,
	dffe17,
	dffe162,
	dffe163,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_0;
input 	sin_o_0;
output 	dffe16;
output 	dffe15;
input 	dffe161;
output 	dffe14;
output 	dffe13;
output 	dffe12;
input 	dffe151;
output 	dffe11;
input 	dffe141;
output 	dffe10;
input 	dffe131;
output 	dffe9;
input 	dffe121;
output 	dffe8;
input 	dffe111;
output 	dffe7;
input 	dffe101;
output 	dffe6;
input 	dffe91;
output 	dffe5;
input 	dffe81;
output 	dffe4;
input 	dffe71;
output 	dffe3;
input 	dffe61;
output 	dffe2;
input 	dffe51;
output 	dffe1;
input 	dffe41;
input 	dffe31;
input 	dffe21;
input 	dffe17;
input 	dffe162;
output 	dffe163;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[15]~q ;
wire \Add0~1_sumout ;
wire \a[14]~q ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \a[13]~q ;
wire \xordvalue[10]~q ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \a[12]~q ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \a[11]~q ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \a[10]~q ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \a[9]~q ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \a[8]~q ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \a[7]~q ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \a[6]~q ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \a[5]~q ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \a[4]~q ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \a[3]~q ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~51 ;
wire \a[2]~q ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~55 ;
wire \a[1]~q ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~59 ;
wire \a[0]~q ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~63 ;


nco_test_lpm_add_sub_51 u0(
	.a_0(a_0),
	.a_15(\a[15]~q ),
	.a_14(\a[14]~q ),
	.a_13(\a[13]~q ),
	.xordvalue_10(\xordvalue[10]~q ),
	.a_12(\a[12]~q ),
	.a_11(\a[11]~q ),
	.a_10(\a[10]~q ),
	.a_9(\a[9]~q ),
	.a_8(\a[8]~q ),
	.a_7(\a[7]~q ),
	.a_6(\a[6]~q ),
	.a_5(\a[5]~q ),
	.a_4(\a[4]~q ),
	.a_3(\a[3]~q ),
	.a_2(\a[2]~q ),
	.a_1(\a[1]~q ),
	.a_01(\a[0]~q ),
	.dffe16(dffe16),
	.dffe15(dffe15),
	.dffe14(dffe14),
	.dffe13(dffe13),
	.dffe12(dffe12),
	.dffe11(dffe11),
	.dffe10(dffe10),
	.dffe9(dffe9),
	.dffe8(dffe8),
	.dffe7(dffe7),
	.dffe6(dffe6),
	.dffe5(dffe5),
	.dffe4(dffe4),
	.dffe3(dffe3),
	.dffe2(dffe2),
	.dffe1(dffe1),
	.dffe161(dffe163),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "on";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~5 .shared_arith = "on";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

dffeas \xordvalue[10] (
	.clk(clk),
	.d(dffe162),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[10]~q ),
	.prn(vcc));
defparam \xordvalue[10] .is_wysiwyg = "true";
defparam \xordvalue[10] .power_up = "low";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~9 .shared_arith = "on";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~13 .shared_arith = "on";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~17 .shared_arith = "on";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "on";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~25 .shared_arith = "on";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~29 .shared_arith = "on";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~33 .shared_arith = "on";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~37 .shared_arith = "on";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(\Add0~47 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~41 .shared_arith = "on";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(\Add0~51 ),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout(\Add0~47 ));
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~45 .shared_arith = "on";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(\Add0~55 ),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout(\Add0~51 ));
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~49 .shared_arith = "on";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(\Add0~59 ),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout(\Add0~55 ));
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~53 .shared_arith = "on";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(\Add0~63 ),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout(\Add0~59 ));
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~57 .shared_arith = "on";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!dffe17),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout(\Add0~63 ));
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add0~61 .shared_arith = "on";

endmodule

module nco_test_lpm_add_sub_51 (
	a_0,
	a_15,
	a_14,
	a_13,
	xordvalue_10,
	a_12,
	a_11,
	a_10,
	a_9,
	a_8,
	a_7,
	a_6,
	a_5,
	a_4,
	a_3,
	a_2,
	a_1,
	a_01,
	dffe16,
	dffe15,
	dffe14,
	dffe13,
	dffe12,
	dffe11,
	dffe10,
	dffe9,
	dffe8,
	dffe7,
	dffe6,
	dffe5,
	dffe4,
	dffe3,
	dffe2,
	dffe1,
	dffe161,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_0;
input 	a_15;
input 	a_14;
input 	a_13;
input 	xordvalue_10;
input 	a_12;
input 	a_11;
input 	a_10;
input 	a_9;
input 	a_8;
input 	a_7;
input 	a_6;
input 	a_5;
input 	a_4;
input 	a_3;
input 	a_2;
input 	a_1;
input 	a_01;
output 	dffe16;
output 	dffe15;
output 	dffe14;
output 	dffe13;
output 	dffe12;
output 	dffe11;
output 	dffe10;
output 	dffe9;
output 	dffe8;
output 	dffe7;
output 	dffe6;
output 	dffe5;
output 	dffe4;
output 	dffe3;
output 	dffe2;
output 	dffe1;
output 	dffe161;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_add_sub_hdg_15 auto_generated(
	.a_0(a_0),
	.a_15(a_15),
	.a_14(a_14),
	.a_13(a_13),
	.xordvalue_10(xordvalue_10),
	.a_12(a_12),
	.a_11(a_11),
	.a_10(a_10),
	.a_9(a_9),
	.a_8(a_8),
	.a_7(a_7),
	.a_6(a_6),
	.a_5(a_5),
	.a_4(a_4),
	.a_3(a_3),
	.a_2(a_2),
	.a_1(a_1),
	.a_01(a_01),
	.dffe161(dffe16),
	.dffe151(dffe15),
	.dffe141(dffe14),
	.dffe131(dffe13),
	.dffe121(dffe12),
	.dffe111(dffe11),
	.dffe101(dffe10),
	.dffe91(dffe9),
	.dffe81(dffe8),
	.dffe71(dffe7),
	.dffe61(dffe6),
	.dffe51(dffe5),
	.dffe41(dffe4),
	.dffe31(dffe3),
	.dffe21(dffe2),
	.dffe17(dffe1),
	.dffe162(dffe161),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module nco_test_add_sub_hdg_15 (
	a_0,
	a_15,
	a_14,
	a_13,
	xordvalue_10,
	a_12,
	a_11,
	a_10,
	a_9,
	a_8,
	a_7,
	a_6,
	a_5,
	a_4,
	a_3,
	a_2,
	a_1,
	a_01,
	dffe161,
	dffe151,
	dffe141,
	dffe131,
	dffe121,
	dffe111,
	dffe101,
	dffe91,
	dffe81,
	dffe71,
	dffe61,
	dffe51,
	dffe41,
	dffe31,
	dffe21,
	dffe17,
	dffe162,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_0;
input 	a_15;
input 	a_14;
input 	a_13;
input 	xordvalue_10;
input 	a_12;
input 	a_11;
input 	a_10;
input 	a_9;
input 	a_8;
input 	a_7;
input 	a_6;
input 	a_5;
input 	a_4;
input 	a_3;
input 	a_2;
input 	a_1;
input 	a_01;
output 	dffe161;
output 	dffe151;
output 	dffe141;
output 	dffe131;
output 	dffe121;
output 	dffe111;
output 	dffe101;
output 	dffe91;
output 	dffe81;
output 	dffe71;
output 	dffe61;
output 	dffe51;
output 	dffe41;
output 	dffe31;
output 	dffe21;
output 	dffe17;
output 	dffe162;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~COUT ;
wire \add_sub_cella[12]~COUT ;
wire \add_sub_cella[13]~COUT ;
wire \add_sub_cella[14]~COUT ;
wire \add_sub_cella[15]~sumout ;
wire \add_sub_cella[14]~sumout ;
wire \add_sub_cella[13]~sumout ;
wire \add_sub_cella[12]~sumout ;
wire \add_sub_cella[11]~sumout ;
wire \add_sub_cella[10]~sumout ;
wire \add_sub_cella[9]~sumout ;
wire \add_sub_cella[8]~sumout ;
wire \add_sub_cella[7]~sumout ;
wire \add_sub_cella[6]~sumout ;
wire \add_sub_cella[5]~sumout ;
wire \add_sub_cella[4]~sumout ;
wire \add_sub_cella[3]~sumout ;
wire \add_sub_cella[2]~sumout ;
wire \add_sub_cella[1]~sumout ;
wire \add_sub_cella[0]~sumout ;


dffeas dffe16(
	.clk(clock),
	.d(\add_sub_cella[15]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe161),
	.prn(vcc));
defparam dffe16.is_wysiwyg = "true";
defparam dffe16.power_up = "low";

dffeas dffe15(
	.clk(clock),
	.d(\add_sub_cella[14]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe151),
	.prn(vcc));
defparam dffe15.is_wysiwyg = "true";
defparam dffe15.power_up = "low";

dffeas dffe14(
	.clk(clock),
	.d(\add_sub_cella[13]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe141),
	.prn(vcc));
defparam dffe14.is_wysiwyg = "true";
defparam dffe14.power_up = "low";

dffeas dffe13(
	.clk(clock),
	.d(\add_sub_cella[12]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe131),
	.prn(vcc));
defparam dffe13.is_wysiwyg = "true";
defparam dffe13.power_up = "low";

dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe17),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

arriav_lcell_comb \dffe16~_wirecell (
	.dataa(!dffe161),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(dffe162),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffe16~_wirecell .extended_lut = "off";
defparam \dffe16~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dffe16~_wirecell .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_01),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(\add_sub_cella[11]~COUT ),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[12] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(\add_sub_cella[11]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[12]~sumout ),
	.cout(\add_sub_cella[12]~COUT ),
	.shareout());
defparam \add_sub_cella[12] .extended_lut = "off";
defparam \add_sub_cella[12] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[12] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[13] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_10),
	.datag(gnd),
	.cin(\add_sub_cella[12]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[13]~sumout ),
	.cout(\add_sub_cella[13]~COUT ),
	.shareout());
defparam \add_sub_cella[13] .extended_lut = "off";
defparam \add_sub_cella[13] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[13] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[14] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(\add_sub_cella[13]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[14]~sumout ),
	.cout(\add_sub_cella[14]~COUT ),
	.shareout());
defparam \add_sub_cella[14] .extended_lut = "off";
defparam \add_sub_cella[14] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[14] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[15] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!a_0),
	.datag(gnd),
	.cin(\add_sub_cella[14]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[15]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[15] .extended_lut = "off";
defparam \add_sub_cella[15] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[15] .shared_arith = "off";

endmodule

module nco_test_cordic_zxor_1p_lpm_16 (
	sin_o_0,
	dffe16,
	dffe15,
	dffe14,
	dffe161,
	dffe13,
	dffe12,
	dffe151,
	dffe11,
	dffe141,
	dffe10,
	dffe131,
	dffe9,
	dffe121,
	dffe8,
	dffe111,
	dffe7,
	dffe101,
	dffe6,
	dffe91,
	dffe5,
	dffe81,
	dffe4,
	dffe71,
	dffe3,
	dffe61,
	dffe2,
	dffe51,
	dffe1,
	dffe41,
	dffe31,
	dffe21,
	dffe17,
	dffe162,
	dffe163,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	sin_o_0;
output 	dffe16;
output 	dffe15;
output 	dffe14;
input 	dffe161;
output 	dffe13;
output 	dffe12;
input 	dffe151;
output 	dffe11;
input 	dffe141;
output 	dffe10;
input 	dffe131;
output 	dffe9;
input 	dffe121;
output 	dffe8;
input 	dffe111;
output 	dffe7;
input 	dffe101;
output 	dffe6;
input 	dffe91;
output 	dffe5;
input 	dffe81;
output 	dffe4;
input 	dffe71;
output 	dffe3;
input 	dffe61;
output 	dffe2;
input 	dffe51;
output 	dffe1;
input 	dffe41;
input 	dffe31;
input 	dffe21;
input 	dffe17;
input 	dffe162;
output 	dffe163;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \a[15]~q ;
wire \xordvalue[0]~q ;
wire \Add0~1_sumout ;
wire \a[14]~q ;
wire \Add0~5_sumout ;
wire \Add0~6 ;
wire \Add0~7 ;
wire \a[13]~q ;
wire \Add0~9_sumout ;
wire \Add0~10 ;
wire \Add0~11 ;
wire \a[12]~q ;
wire \xordvalue[12]~q ;
wire \Add0~13_sumout ;
wire \Add0~14 ;
wire \Add0~15 ;
wire \a[11]~q ;
wire \Add0~17_sumout ;
wire \Add0~18 ;
wire \Add0~19 ;
wire \a[10]~q ;
wire \Add0~21_sumout ;
wire \Add0~22 ;
wire \Add0~23 ;
wire \a[9]~q ;
wire \Add0~25_sumout ;
wire \Add0~26 ;
wire \Add0~27 ;
wire \a[8]~q ;
wire \Add0~29_sumout ;
wire \Add0~30 ;
wire \Add0~31 ;
wire \a[7]~q ;
wire \Add0~33_sumout ;
wire \Add0~34 ;
wire \Add0~35 ;
wire \a[6]~q ;
wire \Add0~37_sumout ;
wire \Add0~38 ;
wire \Add0~39 ;
wire \a[5]~q ;
wire \Add0~41_sumout ;
wire \Add0~42 ;
wire \Add0~43 ;
wire \a[4]~q ;
wire \Add0~45_sumout ;
wire \Add0~46 ;
wire \Add0~47 ;
wire \a[3]~q ;
wire \Add0~49_sumout ;
wire \Add0~50 ;
wire \Add0~51 ;
wire \a[2]~q ;
wire \Add0~53_sumout ;
wire \Add0~54 ;
wire \Add0~55 ;
wire \a[1]~q ;
wire \Add0~57_sumout ;
wire \Add0~58 ;
wire \Add0~59 ;
wire \a[0]~q ;
wire \Add0~61_sumout ;
wire \Add0~62 ;
wire \Add0~63 ;


nco_test_lpm_add_sub_52 u0(
	.a_15(\a[15]~q ),
	.xordvalue_0(\xordvalue[0]~q ),
	.a_14(\a[14]~q ),
	.a_13(\a[13]~q ),
	.a_12(\a[12]~q ),
	.xordvalue_12(\xordvalue[12]~q ),
	.a_11(\a[11]~q ),
	.a_10(\a[10]~q ),
	.a_9(\a[9]~q ),
	.a_8(\a[8]~q ),
	.a_7(\a[7]~q ),
	.a_6(\a[6]~q ),
	.a_5(\a[5]~q ),
	.a_4(\a[4]~q ),
	.a_3(\a[3]~q ),
	.a_2(\a[2]~q ),
	.a_1(\a[1]~q ),
	.a_0(\a[0]~q ),
	.dffe16(dffe16),
	.dffe15(dffe15),
	.dffe14(dffe14),
	.dffe13(dffe13),
	.dffe12(dffe12),
	.dffe11(dffe11),
	.dffe10(dffe10),
	.dffe9(dffe9),
	.dffe8(dffe8),
	.dffe7(dffe7),
	.dffe6(dffe6),
	.dffe5(dffe5),
	.dffe4(dffe4),
	.dffe3(dffe3),
	.dffe2(dffe2),
	.dffe1(dffe1),
	.dffe161(dffe163),
	.clock(clk),
	.reset_n(reset_n),
	.clken(clken));

dffeas \a[15] (
	.clk(clk),
	.d(\Add0~1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[15]~q ),
	.prn(vcc));
defparam \a[15] .is_wysiwyg = "true";
defparam \a[15] .power_up = "low";

dffeas \xordvalue[0] (
	.clk(clk),
	.d(dffe161),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[0]~q ),
	.prn(vcc));
defparam \xordvalue[0] .is_wysiwyg = "true";
defparam \xordvalue[0] .power_up = "low";

arriav_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~6 ),
	.sharein(\Add0~7 ),
	.combout(),
	.sumout(\Add0~1_sumout ),
	.cout(),
	.shareout());
defparam \Add0~1 .extended_lut = "off";
defparam \Add0~1 .lut_mask = 64'h000000000000FF00;
defparam \Add0~1 .shared_arith = "on";

dffeas \a[14] (
	.clk(clk),
	.d(\Add0~5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[14]~q ),
	.prn(vcc));
defparam \a[14] .is_wysiwyg = "true";
defparam \a[14] .power_up = "low";

arriav_lcell_comb \Add0~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe151),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~10 ),
	.sharein(\Add0~11 ),
	.combout(),
	.sumout(\Add0~5_sumout ),
	.cout(\Add0~6 ),
	.shareout(\Add0~7 ));
defparam \Add0~5 .extended_lut = "off";
defparam \Add0~5 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~5 .shared_arith = "on";

dffeas \a[13] (
	.clk(clk),
	.d(\Add0~9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[13]~q ),
	.prn(vcc));
defparam \a[13] .is_wysiwyg = "true";
defparam \a[13] .power_up = "low";

arriav_lcell_comb \Add0~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe141),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~14 ),
	.sharein(\Add0~15 ),
	.combout(),
	.sumout(\Add0~9_sumout ),
	.cout(\Add0~10 ),
	.shareout(\Add0~11 ));
defparam \Add0~9 .extended_lut = "off";
defparam \Add0~9 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~9 .shared_arith = "on";

dffeas \a[12] (
	.clk(clk),
	.d(\Add0~13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[12]~q ),
	.prn(vcc));
defparam \a[12] .is_wysiwyg = "true";
defparam \a[12] .power_up = "low";

dffeas \xordvalue[12] (
	.clk(clk),
	.d(dffe162),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\xordvalue[12]~q ),
	.prn(vcc));
defparam \xordvalue[12] .is_wysiwyg = "true";
defparam \xordvalue[12] .power_up = "low";

arriav_lcell_comb \Add0~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe131),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~18 ),
	.sharein(\Add0~19 ),
	.combout(),
	.sumout(\Add0~13_sumout ),
	.cout(\Add0~14 ),
	.shareout(\Add0~15 ));
defparam \Add0~13 .extended_lut = "off";
defparam \Add0~13 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~13 .shared_arith = "on";

dffeas \a[11] (
	.clk(clk),
	.d(\Add0~17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[11]~q ),
	.prn(vcc));
defparam \a[11] .is_wysiwyg = "true";
defparam \a[11] .power_up = "low";

arriav_lcell_comb \Add0~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe121),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~22 ),
	.sharein(\Add0~23 ),
	.combout(),
	.sumout(\Add0~17_sumout ),
	.cout(\Add0~18 ),
	.shareout(\Add0~19 ));
defparam \Add0~17 .extended_lut = "off";
defparam \Add0~17 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~17 .shared_arith = "on";

dffeas \a[10] (
	.clk(clk),
	.d(\Add0~21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[10]~q ),
	.prn(vcc));
defparam \a[10] .is_wysiwyg = "true";
defparam \a[10] .power_up = "low";

arriav_lcell_comb \Add0~21 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe111),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~26 ),
	.sharein(\Add0~27 ),
	.combout(),
	.sumout(\Add0~21_sumout ),
	.cout(\Add0~22 ),
	.shareout(\Add0~23 ));
defparam \Add0~21 .extended_lut = "off";
defparam \Add0~21 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~21 .shared_arith = "on";

dffeas \a[9] (
	.clk(clk),
	.d(\Add0~25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[9]~q ),
	.prn(vcc));
defparam \a[9] .is_wysiwyg = "true";
defparam \a[9] .power_up = "low";

arriav_lcell_comb \Add0~25 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe101),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~30 ),
	.sharein(\Add0~31 ),
	.combout(),
	.sumout(\Add0~25_sumout ),
	.cout(\Add0~26 ),
	.shareout(\Add0~27 ));
defparam \Add0~25 .extended_lut = "off";
defparam \Add0~25 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~25 .shared_arith = "on";

dffeas \a[8] (
	.clk(clk),
	.d(\Add0~29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[8]~q ),
	.prn(vcc));
defparam \a[8] .is_wysiwyg = "true";
defparam \a[8] .power_up = "low";

arriav_lcell_comb \Add0~29 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe91),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~34 ),
	.sharein(\Add0~35 ),
	.combout(),
	.sumout(\Add0~29_sumout ),
	.cout(\Add0~30 ),
	.shareout(\Add0~31 ));
defparam \Add0~29 .extended_lut = "off";
defparam \Add0~29 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~29 .shared_arith = "on";

dffeas \a[7] (
	.clk(clk),
	.d(\Add0~33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[7]~q ),
	.prn(vcc));
defparam \a[7] .is_wysiwyg = "true";
defparam \a[7] .power_up = "low";

arriav_lcell_comb \Add0~33 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe81),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~38 ),
	.sharein(\Add0~39 ),
	.combout(),
	.sumout(\Add0~33_sumout ),
	.cout(\Add0~34 ),
	.shareout(\Add0~35 ));
defparam \Add0~33 .extended_lut = "off";
defparam \Add0~33 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~33 .shared_arith = "on";

dffeas \a[6] (
	.clk(clk),
	.d(\Add0~37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[6]~q ),
	.prn(vcc));
defparam \a[6] .is_wysiwyg = "true";
defparam \a[6] .power_up = "low";

arriav_lcell_comb \Add0~37 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe71),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~42 ),
	.sharein(\Add0~43 ),
	.combout(),
	.sumout(\Add0~37_sumout ),
	.cout(\Add0~38 ),
	.shareout(\Add0~39 ));
defparam \Add0~37 .extended_lut = "off";
defparam \Add0~37 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~37 .shared_arith = "on";

dffeas \a[5] (
	.clk(clk),
	.d(\Add0~41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[5]~q ),
	.prn(vcc));
defparam \a[5] .is_wysiwyg = "true";
defparam \a[5] .power_up = "low";

arriav_lcell_comb \Add0~41 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe61),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~46 ),
	.sharein(\Add0~47 ),
	.combout(),
	.sumout(\Add0~41_sumout ),
	.cout(\Add0~42 ),
	.shareout(\Add0~43 ));
defparam \Add0~41 .extended_lut = "off";
defparam \Add0~41 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~41 .shared_arith = "on";

dffeas \a[4] (
	.clk(clk),
	.d(\Add0~45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[4]~q ),
	.prn(vcc));
defparam \a[4] .is_wysiwyg = "true";
defparam \a[4] .power_up = "low";

arriav_lcell_comb \Add0~45 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe51),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~50 ),
	.sharein(\Add0~51 ),
	.combout(),
	.sumout(\Add0~45_sumout ),
	.cout(\Add0~46 ),
	.shareout(\Add0~47 ));
defparam \Add0~45 .extended_lut = "off";
defparam \Add0~45 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~45 .shared_arith = "on";

dffeas \a[3] (
	.clk(clk),
	.d(\Add0~49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[3]~q ),
	.prn(vcc));
defparam \a[3] .is_wysiwyg = "true";
defparam \a[3] .power_up = "low";

arriav_lcell_comb \Add0~49 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe41),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~54 ),
	.sharein(\Add0~55 ),
	.combout(),
	.sumout(\Add0~49_sumout ),
	.cout(\Add0~50 ),
	.shareout(\Add0~51 ));
defparam \Add0~49 .extended_lut = "off";
defparam \Add0~49 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~49 .shared_arith = "on";

dffeas \a[2] (
	.clk(clk),
	.d(\Add0~53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[2]~q ),
	.prn(vcc));
defparam \a[2] .is_wysiwyg = "true";
defparam \a[2] .power_up = "low";

arriav_lcell_comb \Add0~53 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe31),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~58 ),
	.sharein(\Add0~59 ),
	.combout(),
	.sumout(\Add0~53_sumout ),
	.cout(\Add0~54 ),
	.shareout(\Add0~55 ));
defparam \Add0~53 .extended_lut = "off";
defparam \Add0~53 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~53 .shared_arith = "on";

dffeas \a[1] (
	.clk(clk),
	.d(\Add0~57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[1]~q ),
	.prn(vcc));
defparam \a[1] .is_wysiwyg = "true";
defparam \a[1] .power_up = "low";

arriav_lcell_comb \Add0~57 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!dffe21),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(\Add0~62 ),
	.sharein(\Add0~63 ),
	.combout(),
	.sumout(\Add0~57_sumout ),
	.cout(\Add0~58 ),
	.shareout(\Add0~59 ));
defparam \Add0~57 .extended_lut = "off";
defparam \Add0~57 .lut_mask = 64'h000000FF0000FF00;
defparam \Add0~57 .shared_arith = "on";

dffeas \a[0] (
	.clk(clk),
	.d(\Add0~61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_0),
	.q(\a[0]~q ),
	.prn(vcc));
defparam \a[0] .is_wysiwyg = "true";
defparam \a[0] .power_up = "low";

arriav_lcell_comb \Add0~61 (
	.dataa(gnd),
	.datab(gnd),
	.datac(!dffe17),
	.datad(!dffe161),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(\Add0~61_sumout ),
	.cout(\Add0~62 ),
	.shareout(\Add0~63 ));
defparam \Add0~61 .extended_lut = "off";
defparam \Add0~61 .lut_mask = 64'h0000FF0F00000FF0;
defparam \Add0~61 .shared_arith = "on";

endmodule

module nco_test_lpm_add_sub_52 (
	a_15,
	xordvalue_0,
	a_14,
	a_13,
	a_12,
	xordvalue_12,
	a_11,
	a_10,
	a_9,
	a_8,
	a_7,
	a_6,
	a_5,
	a_4,
	a_3,
	a_2,
	a_1,
	a_0,
	dffe16,
	dffe15,
	dffe14,
	dffe13,
	dffe12,
	dffe11,
	dffe10,
	dffe9,
	dffe8,
	dffe7,
	dffe6,
	dffe5,
	dffe4,
	dffe3,
	dffe2,
	dffe1,
	dffe161,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_15;
input 	xordvalue_0;
input 	a_14;
input 	a_13;
input 	a_12;
input 	xordvalue_12;
input 	a_11;
input 	a_10;
input 	a_9;
input 	a_8;
input 	a_7;
input 	a_6;
input 	a_5;
input 	a_4;
input 	a_3;
input 	a_2;
input 	a_1;
input 	a_0;
output 	dffe16;
output 	dffe15;
output 	dffe14;
output 	dffe13;
output 	dffe12;
output 	dffe11;
output 	dffe10;
output 	dffe9;
output 	dffe8;
output 	dffe7;
output 	dffe6;
output 	dffe5;
output 	dffe4;
output 	dffe3;
output 	dffe2;
output 	dffe1;
output 	dffe161;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



nco_test_add_sub_hdg_16 auto_generated(
	.a_15(a_15),
	.xordvalue_0(xordvalue_0),
	.a_14(a_14),
	.a_13(a_13),
	.a_12(a_12),
	.xordvalue_12(xordvalue_12),
	.a_11(a_11),
	.a_10(a_10),
	.a_9(a_9),
	.a_8(a_8),
	.a_7(a_7),
	.a_6(a_6),
	.a_5(a_5),
	.a_4(a_4),
	.a_3(a_3),
	.a_2(a_2),
	.a_1(a_1),
	.a_0(a_0),
	.dffe161(dffe16),
	.dffe151(dffe15),
	.dffe141(dffe14),
	.dffe131(dffe13),
	.dffe121(dffe12),
	.dffe111(dffe11),
	.dffe101(dffe10),
	.dffe91(dffe9),
	.dffe81(dffe8),
	.dffe71(dffe7),
	.dffe61(dffe6),
	.dffe51(dffe5),
	.dffe41(dffe4),
	.dffe31(dffe3),
	.dffe21(dffe2),
	.dffe17(dffe1),
	.dffe162(dffe161),
	.clock(clock),
	.reset_n(reset_n),
	.clken(clken));

endmodule

module nco_test_add_sub_hdg_16 (
	a_15,
	xordvalue_0,
	a_14,
	a_13,
	a_12,
	xordvalue_12,
	a_11,
	a_10,
	a_9,
	a_8,
	a_7,
	a_6,
	a_5,
	a_4,
	a_3,
	a_2,
	a_1,
	a_0,
	dffe161,
	dffe151,
	dffe141,
	dffe131,
	dffe121,
	dffe111,
	dffe101,
	dffe91,
	dffe81,
	dffe71,
	dffe61,
	dffe51,
	dffe41,
	dffe31,
	dffe21,
	dffe17,
	dffe162,
	clock,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
input 	a_15;
input 	xordvalue_0;
input 	a_14;
input 	a_13;
input 	a_12;
input 	xordvalue_12;
input 	a_11;
input 	a_10;
input 	a_9;
input 	a_8;
input 	a_7;
input 	a_6;
input 	a_5;
input 	a_4;
input 	a_3;
input 	a_2;
input 	a_1;
input 	a_0;
output 	dffe161;
output 	dffe151;
output 	dffe141;
output 	dffe131;
output 	dffe121;
output 	dffe111;
output 	dffe101;
output 	dffe91;
output 	dffe81;
output 	dffe71;
output 	dffe61;
output 	dffe51;
output 	dffe41;
output 	dffe31;
output 	dffe21;
output 	dffe17;
output 	dffe162;
input 	clock;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \add_sub_cella[0]~2_cout ;
wire \add_sub_cella[0]~COUT ;
wire \add_sub_cella[1]~COUT ;
wire \add_sub_cella[2]~COUT ;
wire \add_sub_cella[3]~COUT ;
wire \add_sub_cella[4]~COUT ;
wire \add_sub_cella[5]~COUT ;
wire \add_sub_cella[6]~COUT ;
wire \add_sub_cella[7]~COUT ;
wire \add_sub_cella[8]~COUT ;
wire \add_sub_cella[9]~COUT ;
wire \add_sub_cella[10]~COUT ;
wire \add_sub_cella[11]~COUT ;
wire \add_sub_cella[12]~COUT ;
wire \add_sub_cella[13]~COUT ;
wire \add_sub_cella[14]~COUT ;
wire \add_sub_cella[15]~sumout ;
wire \add_sub_cella[14]~sumout ;
wire \add_sub_cella[13]~sumout ;
wire \add_sub_cella[12]~sumout ;
wire \add_sub_cella[11]~sumout ;
wire \add_sub_cella[10]~sumout ;
wire \add_sub_cella[9]~sumout ;
wire \add_sub_cella[8]~sumout ;
wire \add_sub_cella[7]~sumout ;
wire \add_sub_cella[6]~sumout ;
wire \add_sub_cella[5]~sumout ;
wire \add_sub_cella[4]~sumout ;
wire \add_sub_cella[3]~sumout ;
wire \add_sub_cella[2]~sumout ;
wire \add_sub_cella[1]~sumout ;
wire \add_sub_cella[0]~sumout ;


dffeas dffe16(
	.clk(clock),
	.d(\add_sub_cella[15]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe161),
	.prn(vcc));
defparam dffe16.is_wysiwyg = "true";
defparam dffe16.power_up = "low";

dffeas dffe15(
	.clk(clock),
	.d(\add_sub_cella[14]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe151),
	.prn(vcc));
defparam dffe15.is_wysiwyg = "true";
defparam dffe15.power_up = "low";

dffeas dffe14(
	.clk(clock),
	.d(\add_sub_cella[13]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe141),
	.prn(vcc));
defparam dffe14.is_wysiwyg = "true";
defparam dffe14.power_up = "low";

dffeas dffe13(
	.clk(clock),
	.d(\add_sub_cella[12]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe131),
	.prn(vcc));
defparam dffe13.is_wysiwyg = "true";
defparam dffe13.power_up = "low";

dffeas dffe12(
	.clk(clock),
	.d(\add_sub_cella[11]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe121),
	.prn(vcc));
defparam dffe12.is_wysiwyg = "true";
defparam dffe12.power_up = "low";

dffeas dffe11(
	.clk(clock),
	.d(\add_sub_cella[10]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe111),
	.prn(vcc));
defparam dffe11.is_wysiwyg = "true";
defparam dffe11.power_up = "low";

dffeas dffe10(
	.clk(clock),
	.d(\add_sub_cella[9]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe101),
	.prn(vcc));
defparam dffe10.is_wysiwyg = "true";
defparam dffe10.power_up = "low";

dffeas dffe9(
	.clk(clock),
	.d(\add_sub_cella[8]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe91),
	.prn(vcc));
defparam dffe9.is_wysiwyg = "true";
defparam dffe9.power_up = "low";

dffeas dffe8(
	.clk(clock),
	.d(\add_sub_cella[7]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe81),
	.prn(vcc));
defparam dffe8.is_wysiwyg = "true";
defparam dffe8.power_up = "low";

dffeas dffe7(
	.clk(clock),
	.d(\add_sub_cella[6]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe71),
	.prn(vcc));
defparam dffe7.is_wysiwyg = "true";
defparam dffe7.power_up = "low";

dffeas dffe6(
	.clk(clock),
	.d(\add_sub_cella[5]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe61),
	.prn(vcc));
defparam dffe6.is_wysiwyg = "true";
defparam dffe6.power_up = "low";

dffeas dffe5(
	.clk(clock),
	.d(\add_sub_cella[4]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe51),
	.prn(vcc));
defparam dffe5.is_wysiwyg = "true";
defparam dffe5.power_up = "low";

dffeas dffe4(
	.clk(clock),
	.d(\add_sub_cella[3]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe41),
	.prn(vcc));
defparam dffe4.is_wysiwyg = "true";
defparam dffe4.power_up = "low";

dffeas dffe3(
	.clk(clock),
	.d(\add_sub_cella[2]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe31),
	.prn(vcc));
defparam dffe3.is_wysiwyg = "true";
defparam dffe3.power_up = "low";

dffeas dffe2(
	.clk(clock),
	.d(\add_sub_cella[1]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe21),
	.prn(vcc));
defparam dffe2.is_wysiwyg = "true";
defparam dffe2.power_up = "low";

dffeas dffe1(
	.clk(clock),
	.d(\add_sub_cella[0]~sumout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(dffe17),
	.prn(vcc));
defparam dffe1.is_wysiwyg = "true";
defparam dffe1.power_up = "low";

arriav_lcell_comb \dffe16~_wirecell (
	.dataa(!dffe161),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(dffe162),
	.sumout(),
	.cout(),
	.shareout());
defparam \dffe16~_wirecell .extended_lut = "off";
defparam \dffe16~_wirecell .lut_mask = 64'hAAAAAAAAAAAAAAAA;
defparam \dffe16~_wirecell .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[0]~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(\add_sub_cella[0]~2_cout ),
	.shareout());
defparam \add_sub_cella[0]~2 .extended_lut = "off";
defparam \add_sub_cella[0]~2 .lut_mask = 64'h0000000000000000;
defparam \add_sub_cella[0]~2 .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[0] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_0),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[0]~2_cout ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[0]~sumout ),
	.cout(\add_sub_cella[0]~COUT ),
	.shareout());
defparam \add_sub_cella[0] .extended_lut = "off";
defparam \add_sub_cella[0] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[0] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[1] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_1),
	.datae(gnd),
	.dataf(!xordvalue_12),
	.datag(gnd),
	.cin(\add_sub_cella[0]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[1]~sumout ),
	.cout(\add_sub_cella[1]~COUT ),
	.shareout());
defparam \add_sub_cella[1] .extended_lut = "off";
defparam \add_sub_cella[1] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[1] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[2] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_2),
	.datae(gnd),
	.dataf(!xordvalue_12),
	.datag(gnd),
	.cin(\add_sub_cella[1]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[2]~sumout ),
	.cout(\add_sub_cella[2]~COUT ),
	.shareout());
defparam \add_sub_cella[2] .extended_lut = "off";
defparam \add_sub_cella[2] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[2] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[3] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_3),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[2]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[3]~sumout ),
	.cout(\add_sub_cella[3]~COUT ),
	.shareout());
defparam \add_sub_cella[3] .extended_lut = "off";
defparam \add_sub_cella[3] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[3] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[4] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_4),
	.datae(gnd),
	.dataf(!xordvalue_12),
	.datag(gnd),
	.cin(\add_sub_cella[3]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[4]~sumout ),
	.cout(\add_sub_cella[4]~COUT ),
	.shareout());
defparam \add_sub_cella[4] .extended_lut = "off";
defparam \add_sub_cella[4] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[4] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[5] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_5),
	.datae(gnd),
	.dataf(!xordvalue_12),
	.datag(gnd),
	.cin(\add_sub_cella[4]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[5]~sumout ),
	.cout(\add_sub_cella[5]~COUT ),
	.shareout());
defparam \add_sub_cella[5] .extended_lut = "off";
defparam \add_sub_cella[5] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[5] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[6] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_6),
	.datae(gnd),
	.dataf(!xordvalue_12),
	.datag(gnd),
	.cin(\add_sub_cella[5]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[6]~sumout ),
	.cout(\add_sub_cella[6]~COUT ),
	.shareout());
defparam \add_sub_cella[6] .extended_lut = "off";
defparam \add_sub_cella[6] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[6] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[7] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_7),
	.datae(gnd),
	.dataf(!xordvalue_12),
	.datag(gnd),
	.cin(\add_sub_cella[6]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[7]~sumout ),
	.cout(\add_sub_cella[7]~COUT ),
	.shareout());
defparam \add_sub_cella[7] .extended_lut = "off";
defparam \add_sub_cella[7] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[7] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[8] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_8),
	.datae(gnd),
	.dataf(!xordvalue_12),
	.datag(gnd),
	.cin(\add_sub_cella[7]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[8]~sumout ),
	.cout(\add_sub_cella[8]~COUT ),
	.shareout());
defparam \add_sub_cella[8] .extended_lut = "off";
defparam \add_sub_cella[8] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[8] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[9] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_9),
	.datae(gnd),
	.dataf(!xordvalue_12),
	.datag(gnd),
	.cin(\add_sub_cella[8]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[9]~sumout ),
	.cout(\add_sub_cella[9]~COUT ),
	.shareout());
defparam \add_sub_cella[9] .extended_lut = "off";
defparam \add_sub_cella[9] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[9] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[10] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_10),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[9]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[10]~sumout ),
	.cout(\add_sub_cella[10]~COUT ),
	.shareout());
defparam \add_sub_cella[10] .extended_lut = "off";
defparam \add_sub_cella[10] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[10] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[11] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_11),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[10]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[11]~sumout ),
	.cout(\add_sub_cella[11]~COUT ),
	.shareout());
defparam \add_sub_cella[11] .extended_lut = "off";
defparam \add_sub_cella[11] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[11] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[12] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_12),
	.datae(gnd),
	.dataf(!xordvalue_12),
	.datag(gnd),
	.cin(\add_sub_cella[11]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[12]~sumout ),
	.cout(\add_sub_cella[12]~COUT ),
	.shareout());
defparam \add_sub_cella[12] .extended_lut = "off";
defparam \add_sub_cella[12] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[12] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[13] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_13),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[12]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[13]~sumout ),
	.cout(\add_sub_cella[13]~COUT ),
	.shareout());
defparam \add_sub_cella[13] .extended_lut = "off";
defparam \add_sub_cella[13] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[13] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[14] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_14),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[13]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[14]~sumout ),
	.cout(\add_sub_cella[14]~COUT ),
	.shareout());
defparam \add_sub_cella[14] .extended_lut = "off";
defparam \add_sub_cella[14] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[14] .shared_arith = "off";

arriav_lcell_comb \add_sub_cella[15] (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!a_15),
	.datae(gnd),
	.dataf(!xordvalue_0),
	.datag(gnd),
	.cin(\add_sub_cella[14]~COUT ),
	.sharein(gnd),
	.combout(),
	.sumout(\add_sub_cella[15]~sumout ),
	.cout(),
	.shareout());
defparam \add_sub_cella[15] .extended_lut = "off";
defparam \add_sub_cella[15] .lut_mask = 64'h000000FF000000FF;
defparam \add_sub_cella[15] .shared_arith = "off";

endmodule

module nco_test_dop_reg (
	sin_o_0,
	sin_o_1,
	sin_o_2,
	sin_o_3,
	sin_o_4,
	sin_o_5,
	sin_o_6,
	sin_o_7,
	sin_o_8,
	sin_o_9,
	sin_o_10,
	sin_o_11,
	sin_o_12,
	sin_o_13,
	sin_o_14,
	sin_o_15,
	sin_o_16,
	sin_o_17,
	cos_o_0,
	cos_o_1,
	cos_o_2,
	cos_o_3,
	cos_o_4,
	cos_o_5,
	cos_o_6,
	cos_o_7,
	cos_o_8,
	cos_o_9,
	cos_o_10,
	cos_o_11,
	cos_o_12,
	cos_o_13,
	cos_o_14,
	cos_o_15,
	cos_o_16,
	cos_o_17,
	sin_o_01,
	sin_o_18,
	sin_o_21,
	sin_o_31,
	sin_o_41,
	sin_o_51,
	sin_o_61,
	sin_o_71,
	sin_o_81,
	sin_o_91,
	sin_o_101,
	sin_o_111,
	sin_o_121,
	sin_o_131,
	sin_o_141,
	sin_o_151,
	sin_o_161,
	sin_o_171,
	cos_o_01,
	cos_o_18,
	cos_o_21,
	cos_o_31,
	cos_o_41,
	cos_o_51,
	cos_o_61,
	cos_o_71,
	cos_o_81,
	cos_o_91,
	cos_o_101,
	cos_o_111,
	cos_o_121,
	cos_o_131,
	cos_o_141,
	cos_o_151,
	cos_o_161,
	cos_o_171,
	sin_o_02,
	clk,
	reset_n,
	clken)/* synthesis synthesis_greybox=1 */;
output 	sin_o_0;
output 	sin_o_1;
output 	sin_o_2;
output 	sin_o_3;
output 	sin_o_4;
output 	sin_o_5;
output 	sin_o_6;
output 	sin_o_7;
output 	sin_o_8;
output 	sin_o_9;
output 	sin_o_10;
output 	sin_o_11;
output 	sin_o_12;
output 	sin_o_13;
output 	sin_o_14;
output 	sin_o_15;
output 	sin_o_16;
output 	sin_o_17;
output 	cos_o_0;
output 	cos_o_1;
output 	cos_o_2;
output 	cos_o_3;
output 	cos_o_4;
output 	cos_o_5;
output 	cos_o_6;
output 	cos_o_7;
output 	cos_o_8;
output 	cos_o_9;
output 	cos_o_10;
output 	cos_o_11;
output 	cos_o_12;
output 	cos_o_13;
output 	cos_o_14;
output 	cos_o_15;
output 	cos_o_16;
output 	cos_o_17;
input 	sin_o_01;
input 	sin_o_18;
input 	sin_o_21;
input 	sin_o_31;
input 	sin_o_41;
input 	sin_o_51;
input 	sin_o_61;
input 	sin_o_71;
input 	sin_o_81;
input 	sin_o_91;
input 	sin_o_101;
input 	sin_o_111;
input 	sin_o_121;
input 	sin_o_131;
input 	sin_o_141;
input 	sin_o_151;
input 	sin_o_161;
input 	sin_o_171;
input 	cos_o_01;
input 	cos_o_18;
input 	cos_o_21;
input 	cos_o_31;
input 	cos_o_41;
input 	cos_o_51;
input 	cos_o_61;
input 	cos_o_71;
input 	cos_o_81;
input 	cos_o_91;
input 	cos_o_101;
input 	cos_o_111;
input 	cos_o_121;
input 	cos_o_131;
input 	cos_o_141;
input 	cos_o_151;
input 	cos_o_161;
input 	cos_o_171;
output 	sin_o_02;
input 	clk;
input 	reset_n;
input 	clken;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas \sin_o[0] (
	.clk(clk),
	.d(sin_o_01),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_02),
	.q(sin_o_0),
	.prn(vcc));
defparam \sin_o[0] .is_wysiwyg = "true";
defparam \sin_o[0] .power_up = "low";

dffeas \sin_o[1] (
	.clk(clk),
	.d(sin_o_18),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_02),
	.q(sin_o_1),
	.prn(vcc));
defparam \sin_o[1] .is_wysiwyg = "true";
defparam \sin_o[1] .power_up = "low";

dffeas \sin_o[2] (
	.clk(clk),
	.d(sin_o_21),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_02),
	.q(sin_o_2),
	.prn(vcc));
defparam \sin_o[2] .is_wysiwyg = "true";
defparam \sin_o[2] .power_up = "low";

dffeas \sin_o[3] (
	.clk(clk),
	.d(sin_o_31),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_02),
	.q(sin_o_3),
	.prn(vcc));
defparam \sin_o[3] .is_wysiwyg = "true";
defparam \sin_o[3] .power_up = "low";

dffeas \sin_o[4] (
	.clk(clk),
	.d(sin_o_41),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_02),
	.q(sin_o_4),
	.prn(vcc));
defparam \sin_o[4] .is_wysiwyg = "true";
defparam \sin_o[4] .power_up = "low";

dffeas \sin_o[5] (
	.clk(clk),
	.d(sin_o_51),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_02),
	.q(sin_o_5),
	.prn(vcc));
defparam \sin_o[5] .is_wysiwyg = "true";
defparam \sin_o[5] .power_up = "low";

dffeas \sin_o[6] (
	.clk(clk),
	.d(sin_o_61),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_02),
	.q(sin_o_6),
	.prn(vcc));
defparam \sin_o[6] .is_wysiwyg = "true";
defparam \sin_o[6] .power_up = "low";

dffeas \sin_o[7] (
	.clk(clk),
	.d(sin_o_71),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_02),
	.q(sin_o_7),
	.prn(vcc));
defparam \sin_o[7] .is_wysiwyg = "true";
defparam \sin_o[7] .power_up = "low";

dffeas \sin_o[8] (
	.clk(clk),
	.d(sin_o_81),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_02),
	.q(sin_o_8),
	.prn(vcc));
defparam \sin_o[8] .is_wysiwyg = "true";
defparam \sin_o[8] .power_up = "low";

dffeas \sin_o[9] (
	.clk(clk),
	.d(sin_o_91),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_02),
	.q(sin_o_9),
	.prn(vcc));
defparam \sin_o[9] .is_wysiwyg = "true";
defparam \sin_o[9] .power_up = "low";

dffeas \sin_o[10] (
	.clk(clk),
	.d(sin_o_101),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_02),
	.q(sin_o_10),
	.prn(vcc));
defparam \sin_o[10] .is_wysiwyg = "true";
defparam \sin_o[10] .power_up = "low";

dffeas \sin_o[11] (
	.clk(clk),
	.d(sin_o_111),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_02),
	.q(sin_o_11),
	.prn(vcc));
defparam \sin_o[11] .is_wysiwyg = "true";
defparam \sin_o[11] .power_up = "low";

dffeas \sin_o[12] (
	.clk(clk),
	.d(sin_o_121),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_02),
	.q(sin_o_12),
	.prn(vcc));
defparam \sin_o[12] .is_wysiwyg = "true";
defparam \sin_o[12] .power_up = "low";

dffeas \sin_o[13] (
	.clk(clk),
	.d(sin_o_131),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_02),
	.q(sin_o_13),
	.prn(vcc));
defparam \sin_o[13] .is_wysiwyg = "true";
defparam \sin_o[13] .power_up = "low";

dffeas \sin_o[14] (
	.clk(clk),
	.d(sin_o_141),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_02),
	.q(sin_o_14),
	.prn(vcc));
defparam \sin_o[14] .is_wysiwyg = "true";
defparam \sin_o[14] .power_up = "low";

dffeas \sin_o[15] (
	.clk(clk),
	.d(sin_o_151),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_02),
	.q(sin_o_15),
	.prn(vcc));
defparam \sin_o[15] .is_wysiwyg = "true";
defparam \sin_o[15] .power_up = "low";

dffeas \sin_o[16] (
	.clk(clk),
	.d(sin_o_161),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_02),
	.q(sin_o_16),
	.prn(vcc));
defparam \sin_o[16] .is_wysiwyg = "true";
defparam \sin_o[16] .power_up = "low";

dffeas \sin_o[17] (
	.clk(clk),
	.d(sin_o_171),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_02),
	.q(sin_o_17),
	.prn(vcc));
defparam \sin_o[17] .is_wysiwyg = "true";
defparam \sin_o[17] .power_up = "low";

dffeas \cos_o[0] (
	.clk(clk),
	.d(cos_o_01),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_02),
	.q(cos_o_0),
	.prn(vcc));
defparam \cos_o[0] .is_wysiwyg = "true";
defparam \cos_o[0] .power_up = "low";

dffeas \cos_o[1] (
	.clk(clk),
	.d(cos_o_18),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_02),
	.q(cos_o_1),
	.prn(vcc));
defparam \cos_o[1] .is_wysiwyg = "true";
defparam \cos_o[1] .power_up = "low";

dffeas \cos_o[2] (
	.clk(clk),
	.d(cos_o_21),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_02),
	.q(cos_o_2),
	.prn(vcc));
defparam \cos_o[2] .is_wysiwyg = "true";
defparam \cos_o[2] .power_up = "low";

dffeas \cos_o[3] (
	.clk(clk),
	.d(cos_o_31),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_02),
	.q(cos_o_3),
	.prn(vcc));
defparam \cos_o[3] .is_wysiwyg = "true";
defparam \cos_o[3] .power_up = "low";

dffeas \cos_o[4] (
	.clk(clk),
	.d(cos_o_41),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_02),
	.q(cos_o_4),
	.prn(vcc));
defparam \cos_o[4] .is_wysiwyg = "true";
defparam \cos_o[4] .power_up = "low";

dffeas \cos_o[5] (
	.clk(clk),
	.d(cos_o_51),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_02),
	.q(cos_o_5),
	.prn(vcc));
defparam \cos_o[5] .is_wysiwyg = "true";
defparam \cos_o[5] .power_up = "low";

dffeas \cos_o[6] (
	.clk(clk),
	.d(cos_o_61),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_02),
	.q(cos_o_6),
	.prn(vcc));
defparam \cos_o[6] .is_wysiwyg = "true";
defparam \cos_o[6] .power_up = "low";

dffeas \cos_o[7] (
	.clk(clk),
	.d(cos_o_71),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_02),
	.q(cos_o_7),
	.prn(vcc));
defparam \cos_o[7] .is_wysiwyg = "true";
defparam \cos_o[7] .power_up = "low";

dffeas \cos_o[8] (
	.clk(clk),
	.d(cos_o_81),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_02),
	.q(cos_o_8),
	.prn(vcc));
defparam \cos_o[8] .is_wysiwyg = "true";
defparam \cos_o[8] .power_up = "low";

dffeas \cos_o[9] (
	.clk(clk),
	.d(cos_o_91),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_02),
	.q(cos_o_9),
	.prn(vcc));
defparam \cos_o[9] .is_wysiwyg = "true";
defparam \cos_o[9] .power_up = "low";

dffeas \cos_o[10] (
	.clk(clk),
	.d(cos_o_101),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_02),
	.q(cos_o_10),
	.prn(vcc));
defparam \cos_o[10] .is_wysiwyg = "true";
defparam \cos_o[10] .power_up = "low";

dffeas \cos_o[11] (
	.clk(clk),
	.d(cos_o_111),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_02),
	.q(cos_o_11),
	.prn(vcc));
defparam \cos_o[11] .is_wysiwyg = "true";
defparam \cos_o[11] .power_up = "low";

dffeas \cos_o[12] (
	.clk(clk),
	.d(cos_o_121),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_02),
	.q(cos_o_12),
	.prn(vcc));
defparam \cos_o[12] .is_wysiwyg = "true";
defparam \cos_o[12] .power_up = "low";

dffeas \cos_o[13] (
	.clk(clk),
	.d(cos_o_131),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_02),
	.q(cos_o_13),
	.prn(vcc));
defparam \cos_o[13] .is_wysiwyg = "true";
defparam \cos_o[13] .power_up = "low";

dffeas \cos_o[14] (
	.clk(clk),
	.d(cos_o_141),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_02),
	.q(cos_o_14),
	.prn(vcc));
defparam \cos_o[14] .is_wysiwyg = "true";
defparam \cos_o[14] .power_up = "low";

dffeas \cos_o[15] (
	.clk(clk),
	.d(cos_o_151),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_02),
	.q(cos_o_15),
	.prn(vcc));
defparam \cos_o[15] .is_wysiwyg = "true";
defparam \cos_o[15] .power_up = "low";

dffeas \cos_o[16] (
	.clk(clk),
	.d(cos_o_161),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_02),
	.q(cos_o_16),
	.prn(vcc));
defparam \cos_o[16] .is_wysiwyg = "true";
defparam \cos_o[16] .power_up = "low";

dffeas \cos_o[17] (
	.clk(clk),
	.d(cos_o_171),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(sin_o_02),
	.q(cos_o_17),
	.prn(vcc));
defparam \cos_o[17] .is_wysiwyg = "true";
defparam \cos_o[17] .power_up = "low";

arriav_lcell_comb \sin_o[0]~0 (
	.dataa(!reset_n),
	.datab(!clken),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(sin_o_02),
	.sumout(),
	.cout(),
	.shareout());
defparam \sin_o[0]~0 .extended_lut = "off";
defparam \sin_o[0]~0 .lut_mask = 64'hBBBBBBBBBBBBBBBB;
defparam \sin_o[0]~0 .shared_arith = "off";

endmodule
