
module GBUF_RST (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
