
module mypll (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
